library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4e0c287",
    12 => x"86c0c64e",
    13 => x"49c4e0c2",
    14 => x"48f8cdc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087ffd6",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"d4ff1e4f",
    50 => x"78ffc348",
    51 => x"66c45168",
    52 => x"c888c148",
    53 => x"987058a6",
    54 => x"2687eb05",
    55 => x"1e731e4f",
    56 => x"c34bd4ff",
    57 => x"4a6b7bff",
    58 => x"6b7bffc3",
    59 => x"7232c849",
    60 => x"7bffc3b1",
    61 => x"31c84a6b",
    62 => x"ffc3b271",
    63 => x"c8496b7b",
    64 => x"71b17232",
    65 => x"2687c448",
    66 => x"264c264d",
    67 => x"0e4f264b",
    68 => x"5d5c5b5e",
    69 => x"ff4a710e",
    70 => x"49724cd4",
    71 => x"7199ffc3",
    72 => x"f8cdc27c",
    73 => x"87c805bf",
    74 => x"c94866d0",
    75 => x"58a6d430",
    76 => x"d84966d0",
    77 => x"99ffc329",
    78 => x"66d07c71",
    79 => x"c329d049",
    80 => x"7c7199ff",
    81 => x"c84966d0",
    82 => x"99ffc329",
    83 => x"66d07c71",
    84 => x"99ffc349",
    85 => x"49727c71",
    86 => x"ffc329d0",
    87 => x"6c7c7199",
    88 => x"fff0c94b",
    89 => x"abffc34d",
    90 => x"c387d005",
    91 => x"4b6c7cff",
    92 => x"c6028dc1",
    93 => x"abffc387",
    94 => x"7387f002",
    95 => x"87c7fe48",
    96 => x"ff49c01e",
    97 => x"ffc348d4",
    98 => x"c381c178",
    99 => x"04a9b7c8",
   100 => x"4f2687f1",
   101 => x"e71e731e",
   102 => x"dff8c487",
   103 => x"c01ec04b",
   104 => x"f7c1f0ff",
   105 => x"87e7fd49",
   106 => x"a8c186c4",
   107 => x"87eac005",
   108 => x"c348d4ff",
   109 => x"c0c178ff",
   110 => x"c0c0c0c0",
   111 => x"f0e1c01e",
   112 => x"fd49e9c1",
   113 => x"86c487c9",
   114 => x"ca059870",
   115 => x"48d4ff87",
   116 => x"c178ffc3",
   117 => x"fe87cb48",
   118 => x"8bc187e6",
   119 => x"87fdfe05",
   120 => x"e6fc48c0",
   121 => x"1e731e87",
   122 => x"c348d4ff",
   123 => x"4bd378ff",
   124 => x"ffc01ec0",
   125 => x"49c1c1f0",
   126 => x"c487d4fc",
   127 => x"05987086",
   128 => x"d4ff87ca",
   129 => x"78ffc348",
   130 => x"87cb48c1",
   131 => x"c187f1fd",
   132 => x"dbff058b",
   133 => x"fb48c087",
   134 => x"5e0e87f1",
   135 => x"ff0e5c5b",
   136 => x"dbfd4cd4",
   137 => x"1eeac687",
   138 => x"c1f0e1c0",
   139 => x"defb49c8",
   140 => x"c186c487",
   141 => x"87c802a8",
   142 => x"c087eafe",
   143 => x"87e2c148",
   144 => x"7087dafa",
   145 => x"ffffcf49",
   146 => x"a9eac699",
   147 => x"fe87c802",
   148 => x"48c087d3",
   149 => x"c387cbc1",
   150 => x"f1c07cff",
   151 => x"87f4fc4b",
   152 => x"c0029870",
   153 => x"1ec087eb",
   154 => x"c1f0ffc0",
   155 => x"defa49fa",
   156 => x"7086c487",
   157 => x"87d90598",
   158 => x"6c7cffc3",
   159 => x"7cffc349",
   160 => x"c17c7c7c",
   161 => x"c40299c0",
   162 => x"d548c187",
   163 => x"d148c087",
   164 => x"05abc287",
   165 => x"48c087c4",
   166 => x"8bc187c8",
   167 => x"87fdfe05",
   168 => x"e4f948c0",
   169 => x"1e731e87",
   170 => x"48f8cdc2",
   171 => x"4bc778c1",
   172 => x"c248d0ff",
   173 => x"87c8fb78",
   174 => x"c348d0ff",
   175 => x"c01ec078",
   176 => x"c0c1d0e5",
   177 => x"87c7f949",
   178 => x"a8c186c4",
   179 => x"4b87c105",
   180 => x"c505abc2",
   181 => x"c048c087",
   182 => x"8bc187f9",
   183 => x"87d0ff05",
   184 => x"c287f7fc",
   185 => x"7058fccd",
   186 => x"87cd0598",
   187 => x"ffc01ec1",
   188 => x"49d0c1f0",
   189 => x"c487d8f8",
   190 => x"48d4ff86",
   191 => x"c278ffc3",
   192 => x"cec287fe",
   193 => x"d0ff58c0",
   194 => x"ff78c248",
   195 => x"ffc348d4",
   196 => x"f748c178",
   197 => x"ff1e87f5",
   198 => x"d0ff4ad4",
   199 => x"78d1c448",
   200 => x"c17affc3",
   201 => x"87f80589",
   202 => x"731e4f26",
   203 => x"c54b711e",
   204 => x"4adfcdee",
   205 => x"c348d4ff",
   206 => x"486878ff",
   207 => x"02a8fec3",
   208 => x"8ac187c5",
   209 => x"7287ed05",
   210 => x"87c5059a",
   211 => x"eac048c0",
   212 => x"029b7387",
   213 => x"66c887cc",
   214 => x"f549731e",
   215 => x"86c487e7",
   216 => x"66c887c6",
   217 => x"87eefe49",
   218 => x"c348d4ff",
   219 => x"737878ff",
   220 => x"87c5059b",
   221 => x"d048d0ff",
   222 => x"f648c178",
   223 => x"731e87cd",
   224 => x"c04a711e",
   225 => x"48d4ff4b",
   226 => x"ff78ffc3",
   227 => x"c3c448d0",
   228 => x"48d4ff78",
   229 => x"7278ffc3",
   230 => x"f0ffc01e",
   231 => x"f549d1c1",
   232 => x"86c487ed",
   233 => x"cd059870",
   234 => x"1ec0c887",
   235 => x"fd4966cc",
   236 => x"86c487f8",
   237 => x"d0ff4b70",
   238 => x"7378c248",
   239 => x"87cbf548",
   240 => x"5c5b5e0e",
   241 => x"1ec00e5d",
   242 => x"c1f0ffc0",
   243 => x"fef449c9",
   244 => x"c21ed287",
   245 => x"fd49c0ce",
   246 => x"86c887d0",
   247 => x"84c14cc0",
   248 => x"04acb7d2",
   249 => x"cec287f8",
   250 => x"49bf97c0",
   251 => x"c199c0c3",
   252 => x"c005a9c0",
   253 => x"cec287e7",
   254 => x"49bf97c7",
   255 => x"cec231d0",
   256 => x"4abf97c8",
   257 => x"b17232c8",
   258 => x"97c9cec2",
   259 => x"71b14abf",
   260 => x"ffffcf4c",
   261 => x"84c19cff",
   262 => x"e7c134ca",
   263 => x"c9cec287",
   264 => x"c149bf97",
   265 => x"c299c631",
   266 => x"bf97cace",
   267 => x"2ab7c74a",
   268 => x"cec2b172",
   269 => x"4abf97c5",
   270 => x"c29dcf4d",
   271 => x"bf97c6ce",
   272 => x"ca9ac34a",
   273 => x"c7cec232",
   274 => x"c24bbf97",
   275 => x"c2b27333",
   276 => x"bf97c8ce",
   277 => x"9bc0c34b",
   278 => x"732bb7c6",
   279 => x"c181c2b2",
   280 => x"70307148",
   281 => x"7548c149",
   282 => x"724d7030",
   283 => x"7184c14c",
   284 => x"b7c0c894",
   285 => x"87cc06ad",
   286 => x"2db734c1",
   287 => x"adb7c0c8",
   288 => x"87f4ff01",
   289 => x"fef14874",
   290 => x"5b5e0e87",
   291 => x"f80e5d5c",
   292 => x"e6d6c286",
   293 => x"c278c048",
   294 => x"c01edece",
   295 => x"87defb49",
   296 => x"987086c4",
   297 => x"c087c505",
   298 => x"87cec948",
   299 => x"7ec14dc0",
   300 => x"bfe9edc0",
   301 => x"d4cfc249",
   302 => x"4bc8714a",
   303 => x"7087ebee",
   304 => x"87c20598",
   305 => x"edc07ec0",
   306 => x"c249bfe5",
   307 => x"714af0cf",
   308 => x"d5ee4bc8",
   309 => x"05987087",
   310 => x"7ec087c2",
   311 => x"fdc0026e",
   312 => x"e4d5c287",
   313 => x"d6c24dbf",
   314 => x"7ebf9fdc",
   315 => x"ead6c548",
   316 => x"87c705a8",
   317 => x"bfe4d5c2",
   318 => x"6e87ce4d",
   319 => x"d5e9ca48",
   320 => x"87c502a8",
   321 => x"f1c748c0",
   322 => x"decec287",
   323 => x"f949751e",
   324 => x"86c487ec",
   325 => x"c5059870",
   326 => x"c748c087",
   327 => x"edc087dc",
   328 => x"c249bfe5",
   329 => x"714af0cf",
   330 => x"fdec4bc8",
   331 => x"05987087",
   332 => x"d6c287c8",
   333 => x"78c148e6",
   334 => x"edc087da",
   335 => x"c249bfe9",
   336 => x"714ad4cf",
   337 => x"e1ec4bc8",
   338 => x"02987087",
   339 => x"c087c5c0",
   340 => x"87e6c648",
   341 => x"97dcd6c2",
   342 => x"d5c149bf",
   343 => x"cdc005a9",
   344 => x"ddd6c287",
   345 => x"c249bf97",
   346 => x"c002a9ea",
   347 => x"48c087c5",
   348 => x"c287c7c6",
   349 => x"bf97dece",
   350 => x"e9c3487e",
   351 => x"cec002a8",
   352 => x"c3486e87",
   353 => x"c002a8eb",
   354 => x"48c087c5",
   355 => x"c287ebc5",
   356 => x"bf97e9ce",
   357 => x"c0059949",
   358 => x"cec287cc",
   359 => x"49bf97ea",
   360 => x"c002a9c2",
   361 => x"48c087c5",
   362 => x"c287cfc5",
   363 => x"bf97ebce",
   364 => x"e2d6c248",
   365 => x"484c7058",
   366 => x"d6c288c1",
   367 => x"cec258e6",
   368 => x"49bf97ec",
   369 => x"cec28175",
   370 => x"4abf97ed",
   371 => x"a17232c8",
   372 => x"f3dac27e",
   373 => x"c2786e48",
   374 => x"bf97eece",
   375 => x"58a6c848",
   376 => x"bfe6d6c2",
   377 => x"87d4c202",
   378 => x"bfe5edc0",
   379 => x"f0cfc249",
   380 => x"4bc8714a",
   381 => x"7087f3e9",
   382 => x"c5c00298",
   383 => x"c348c087",
   384 => x"d6c287f8",
   385 => x"c24cbfde",
   386 => x"c25cc7db",
   387 => x"bf97c3cf",
   388 => x"c231c849",
   389 => x"bf97c2cf",
   390 => x"c249a14a",
   391 => x"bf97c4cf",
   392 => x"7232d04a",
   393 => x"cfc249a1",
   394 => x"4abf97c5",
   395 => x"a17232d8",
   396 => x"9166c449",
   397 => x"bff3dac2",
   398 => x"fbdac281",
   399 => x"cbcfc259",
   400 => x"c84abf97",
   401 => x"cacfc232",
   402 => x"a24bbf97",
   403 => x"cccfc24a",
   404 => x"d04bbf97",
   405 => x"4aa27333",
   406 => x"97cdcfc2",
   407 => x"9bcf4bbf",
   408 => x"a27333d8",
   409 => x"ffdac24a",
   410 => x"fbdac25a",
   411 => x"8ac24abf",
   412 => x"dac29274",
   413 => x"a17248ff",
   414 => x"87cac178",
   415 => x"97f0cec2",
   416 => x"31c849bf",
   417 => x"97efcec2",
   418 => x"49a14abf",
   419 => x"59eed6c2",
   420 => x"bfead6c2",
   421 => x"c731c549",
   422 => x"29c981ff",
   423 => x"59c7dbc2",
   424 => x"97f5cec2",
   425 => x"32c84abf",
   426 => x"97f4cec2",
   427 => x"4aa24bbf",
   428 => x"6e9266c4",
   429 => x"c3dbc282",
   430 => x"fbdac25a",
   431 => x"c278c048",
   432 => x"7248f7da",
   433 => x"dbc278a1",
   434 => x"dac248c7",
   435 => x"c278bffb",
   436 => x"c248cbdb",
   437 => x"78bfffda",
   438 => x"bfe6d6c2",
   439 => x"87c9c002",
   440 => x"30c44874",
   441 => x"c9c07e70",
   442 => x"c3dbc287",
   443 => x"30c448bf",
   444 => x"d6c27e70",
   445 => x"786e48ea",
   446 => x"8ef848c1",
   447 => x"4c264d26",
   448 => x"4f264b26",
   449 => x"5c5b5e0e",
   450 => x"4a710e5d",
   451 => x"bfe6d6c2",
   452 => x"7287cb02",
   453 => x"722bc74b",
   454 => x"9cffc14c",
   455 => x"4b7287c9",
   456 => x"4c722bc8",
   457 => x"c29cffc3",
   458 => x"83bff3da",
   459 => x"bfe1edc0",
   460 => x"87d902ab",
   461 => x"5be5edc0",
   462 => x"1edecec2",
   463 => x"fdf04973",
   464 => x"7086c487",
   465 => x"87c50598",
   466 => x"e6c048c0",
   467 => x"e6d6c287",
   468 => x"87d202bf",
   469 => x"91c44974",
   470 => x"81decec2",
   471 => x"ffcf4d69",
   472 => x"9dffffff",
   473 => x"497487cb",
   474 => x"cec291c2",
   475 => x"699f81de",
   476 => x"fe48754d",
   477 => x"5e0e87c6",
   478 => x"0e5d5c5b",
   479 => x"c04d711e",
   480 => x"c849c11e",
   481 => x"86c487c4",
   482 => x"029c4c70",
   483 => x"c287c0c1",
   484 => x"754aeed6",
   485 => x"87f7e249",
   486 => x"c0029870",
   487 => x"4a7487f1",
   488 => x"4bcb4975",
   489 => x"7087dde3",
   490 => x"e2c00298",
   491 => x"741ec087",
   492 => x"87c7029c",
   493 => x"c048a6c4",
   494 => x"c487c578",
   495 => x"78c148a6",
   496 => x"c74966c4",
   497 => x"86c487c4",
   498 => x"059c4c70",
   499 => x"7487c0ff",
   500 => x"e7fc2648",
   501 => x"5b5e0e87",
   502 => x"1e0e5d5c",
   503 => x"059b4b71",
   504 => x"48c087c5",
   505 => x"c887e5c1",
   506 => x"7dc04da3",
   507 => x"c70266d4",
   508 => x"9766d487",
   509 => x"87c505bf",
   510 => x"cfc148c0",
   511 => x"4966d487",
   512 => x"7087f3fd",
   513 => x"c1029c4c",
   514 => x"a4dc87c0",
   515 => x"da7d6949",
   516 => x"a3c449a4",
   517 => x"7a699f4a",
   518 => x"bfe6d6c2",
   519 => x"d487d202",
   520 => x"699f49a4",
   521 => x"ffffc049",
   522 => x"d0487199",
   523 => x"c27e7030",
   524 => x"6e7ec087",
   525 => x"806a4849",
   526 => x"7bc07a70",
   527 => x"6a49a3cc",
   528 => x"49a3d079",
   529 => x"487479c0",
   530 => x"48c087c2",
   531 => x"87ecfa26",
   532 => x"5c5b5e0e",
   533 => x"4c710e5d",
   534 => x"48e1edc0",
   535 => x"9c7478ff",
   536 => x"87cac102",
   537 => x"6949a4c8",
   538 => x"87c2c102",
   539 => x"6c4a66d0",
   540 => x"a6d48249",
   541 => x"4d66d05a",
   542 => x"e2d6c2b9",
   543 => x"baff4abf",
   544 => x"99719972",
   545 => x"87e4c002",
   546 => x"6b4ba4c4",
   547 => x"87f4f949",
   548 => x"d6c27b70",
   549 => x"6c49bfde",
   550 => x"757c7181",
   551 => x"e2d6c2b9",
   552 => x"baff4abf",
   553 => x"99719972",
   554 => x"87dcff05",
   555 => x"cbf97c75",
   556 => x"1e731e87",
   557 => x"029b4b71",
   558 => x"a3c887c7",
   559 => x"c5056949",
   560 => x"c048c087",
   561 => x"dac287eb",
   562 => x"c44abff7",
   563 => x"496949a3",
   564 => x"d6c289c2",
   565 => x"7191bfde",
   566 => x"d6c24aa2",
   567 => x"6b49bfe2",
   568 => x"4aa27199",
   569 => x"721e66c8",
   570 => x"87d2ea49",
   571 => x"497086c4",
   572 => x"87ccf848",
   573 => x"711e731e",
   574 => x"c0029b4b",
   575 => x"dbc287e4",
   576 => x"4a735bcb",
   577 => x"d6c28ac2",
   578 => x"9249bfde",
   579 => x"bff7dac2",
   580 => x"c2807248",
   581 => x"7158cfdb",
   582 => x"c230c448",
   583 => x"c058eed6",
   584 => x"dbc287ed",
   585 => x"dac248c7",
   586 => x"c278bffb",
   587 => x"c248cbdb",
   588 => x"78bfffda",
   589 => x"bfe6d6c2",
   590 => x"c287c902",
   591 => x"49bfded6",
   592 => x"87c731c4",
   593 => x"bfc3dbc2",
   594 => x"c231c449",
   595 => x"f659eed6",
   596 => x"5e0e87ee",
   597 => x"710e5c5b",
   598 => x"724bc04a",
   599 => x"e1c0029a",
   600 => x"49a2da87",
   601 => x"c24b699f",
   602 => x"02bfe6d6",
   603 => x"a2d487cf",
   604 => x"49699f49",
   605 => x"ffffc04c",
   606 => x"c234d09c",
   607 => x"744cc087",
   608 => x"4973b349",
   609 => x"f587edfd",
   610 => x"5e0e87f4",
   611 => x"0e5d5c5b",
   612 => x"4a7186f4",
   613 => x"9a727ec0",
   614 => x"c287d802",
   615 => x"c048dace",
   616 => x"d2cec278",
   617 => x"cbdbc248",
   618 => x"cec278bf",
   619 => x"dbc248d6",
   620 => x"c278bfc7",
   621 => x"c048fbd6",
   622 => x"ead6c250",
   623 => x"cec249bf",
   624 => x"714abfda",
   625 => x"ffc303aa",
   626 => x"cf497287",
   627 => x"e0c00599",
   628 => x"decec287",
   629 => x"d2cec21e",
   630 => x"cec249bf",
   631 => x"a1c148d2",
   632 => x"d9e67178",
   633 => x"c086c487",
   634 => x"c248dded",
   635 => x"cc78dece",
   636 => x"ddedc087",
   637 => x"e0c048bf",
   638 => x"e1edc080",
   639 => x"dacec258",
   640 => x"80c148bf",
   641 => x"58decec2",
   642 => x"000b5d27",
   643 => x"bf97bf00",
   644 => x"c2029d4d",
   645 => x"e5c387e2",
   646 => x"dbc202ad",
   647 => x"ddedc087",
   648 => x"a3cb4bbf",
   649 => x"cf4c1149",
   650 => x"d2c105ac",
   651 => x"df497587",
   652 => x"cd89c199",
   653 => x"eed6c291",
   654 => x"4aa3c181",
   655 => x"a3c35112",
   656 => x"c551124a",
   657 => x"51124aa3",
   658 => x"124aa3c7",
   659 => x"4aa3c951",
   660 => x"a3ce5112",
   661 => x"d051124a",
   662 => x"51124aa3",
   663 => x"124aa3d2",
   664 => x"4aa3d451",
   665 => x"a3d65112",
   666 => x"d851124a",
   667 => x"51124aa3",
   668 => x"124aa3dc",
   669 => x"4aa3de51",
   670 => x"7ec15112",
   671 => x"7487f9c0",
   672 => x"0599c849",
   673 => x"7487eac0",
   674 => x"0599d049",
   675 => x"66dc87d0",
   676 => x"87cac002",
   677 => x"66dc4973",
   678 => x"0298700f",
   679 => x"056e87d3",
   680 => x"c287c6c0",
   681 => x"c048eed6",
   682 => x"ddedc050",
   683 => x"e7c248bf",
   684 => x"fbd6c287",
   685 => x"7e50c048",
   686 => x"bfead6c2",
   687 => x"dacec249",
   688 => x"aa714abf",
   689 => x"87c1fc04",
   690 => x"bfcbdbc2",
   691 => x"87c8c005",
   692 => x"bfe6d6c2",
   693 => x"87fec102",
   694 => x"48e1edc0",
   695 => x"cec278ff",
   696 => x"f049bfd6",
   697 => x"497087de",
   698 => x"59dacec2",
   699 => x"c248a6c4",
   700 => x"78bfd6ce",
   701 => x"bfe6d6c2",
   702 => x"87d8c002",
   703 => x"cf4966c4",
   704 => x"f8ffffff",
   705 => x"c002a999",
   706 => x"4dc087c5",
   707 => x"c187e1c0",
   708 => x"87dcc04d",
   709 => x"cf4966c4",
   710 => x"a999f8ff",
   711 => x"87c8c002",
   712 => x"c048a6c8",
   713 => x"87c5c078",
   714 => x"c148a6c8",
   715 => x"4d66c878",
   716 => x"c0059d75",
   717 => x"66c487e0",
   718 => x"c289c249",
   719 => x"4abfded6",
   720 => x"f7dac291",
   721 => x"cec24abf",
   722 => x"a17248d2",
   723 => x"dacec278",
   724 => x"f978c048",
   725 => x"48c087e3",
   726 => x"dfee8ef4",
   727 => x"00000087",
   728 => x"ffffff00",
   729 => x"000b6dff",
   730 => x"000b7600",
   731 => x"54414600",
   732 => x"20203233",
   733 => x"41460020",
   734 => x"20363154",
   735 => x"1e002020",
   736 => x"c348d4ff",
   737 => x"486878ff",
   738 => x"ff1e4f26",
   739 => x"ffc348d4",
   740 => x"48d0ff78",
   741 => x"ff78e1c8",
   742 => x"78d448d4",
   743 => x"48cfdbc2",
   744 => x"50bfd4ff",
   745 => x"ff1e4f26",
   746 => x"e0c048d0",
   747 => x"1e4f2678",
   748 => x"7087ccff",
   749 => x"c6029949",
   750 => x"a9fbc087",
   751 => x"7187f105",
   752 => x"0e4f2648",
   753 => x"0e5c5b5e",
   754 => x"4cc04b71",
   755 => x"7087f0fe",
   756 => x"c0029949",
   757 => x"ecc087f9",
   758 => x"f2c002a9",
   759 => x"a9fbc087",
   760 => x"87ebc002",
   761 => x"acb766cc",
   762 => x"d087c703",
   763 => x"87c20266",
   764 => x"99715371",
   765 => x"c187c202",
   766 => x"87c3fe84",
   767 => x"02994970",
   768 => x"ecc087cd",
   769 => x"87c702a9",
   770 => x"05a9fbc0",
   771 => x"d087d5ff",
   772 => x"87c30266",
   773 => x"c07b97c0",
   774 => x"c405a9ec",
   775 => x"c54a7487",
   776 => x"c04a7487",
   777 => x"48728a0a",
   778 => x"4d2687c2",
   779 => x"4b264c26",
   780 => x"fd1e4f26",
   781 => x"497087c9",
   782 => x"a9b7f0c0",
   783 => x"c087ca04",
   784 => x"01a9b7f9",
   785 => x"f0c087c3",
   786 => x"b7c1c189",
   787 => x"87ca04a9",
   788 => x"a9b7dac1",
   789 => x"c087c301",
   790 => x"487189f7",
   791 => x"5e0e4f26",
   792 => x"710e5c5b",
   793 => x"4cd4ff4a",
   794 => x"eac04972",
   795 => x"9b4b7087",
   796 => x"c187c202",
   797 => x"48d0ff8b",
   798 => x"c178c5c8",
   799 => x"49737cd5",
   800 => x"cdc231c6",
   801 => x"4abf97ca",
   802 => x"70b07148",
   803 => x"48d0ff7c",
   804 => x"487378c4",
   805 => x"0e87d5fe",
   806 => x"5d5c5b5e",
   807 => x"7186f80e",
   808 => x"fb7ec04c",
   809 => x"4bc087e4",
   810 => x"97c4f5c0",
   811 => x"a9c049bf",
   812 => x"fb87cf04",
   813 => x"83c187f9",
   814 => x"97c4f5c0",
   815 => x"06ab49bf",
   816 => x"f5c087f1",
   817 => x"02bf97c4",
   818 => x"f2fa87cf",
   819 => x"99497087",
   820 => x"c087c602",
   821 => x"f105a9ec",
   822 => x"fa4bc087",
   823 => x"4d7087e1",
   824 => x"c887dcfa",
   825 => x"d6fa58a6",
   826 => x"c14a7087",
   827 => x"49a4c883",
   828 => x"ad496997",
   829 => x"c087c702",
   830 => x"c005adff",
   831 => x"a4c987e7",
   832 => x"49699749",
   833 => x"02a966c4",
   834 => x"c04887c7",
   835 => x"d405a8ff",
   836 => x"49a4ca87",
   837 => x"aa496997",
   838 => x"c087c602",
   839 => x"c405aaff",
   840 => x"d07ec187",
   841 => x"adecc087",
   842 => x"c087c602",
   843 => x"c405adfb",
   844 => x"c14bc087",
   845 => x"fe026e7e",
   846 => x"e9f987e1",
   847 => x"f8487387",
   848 => x"87e6fb8e",
   849 => x"5b5e0e00",
   850 => x"1e0e5d5c",
   851 => x"4cc04b71",
   852 => x"c004ab4d",
   853 => x"f2c087e8",
   854 => x"9d751ed7",
   855 => x"c087c402",
   856 => x"c187c24a",
   857 => x"f049724a",
   858 => x"86c487e0",
   859 => x"84c17e70",
   860 => x"87c2056e",
   861 => x"85c14c73",
   862 => x"ff06ac73",
   863 => x"486e87d8",
   864 => x"264d2626",
   865 => x"264b264c",
   866 => x"5b5e0e4f",
   867 => x"1e0e5d5c",
   868 => x"de494c71",
   869 => x"e9dbc291",
   870 => x"9785714d",
   871 => x"ddc1026d",
   872 => x"d4dbc287",
   873 => x"82744abf",
   874 => x"d8fe4972",
   875 => x"6e7e7087",
   876 => x"87f3c002",
   877 => x"4bdcdbc2",
   878 => x"49cb4a6e",
   879 => x"87e8cbff",
   880 => x"93cb4b74",
   881 => x"83eed8c1",
   882 => x"f8c083c4",
   883 => x"49747bc2",
   884 => x"87d8c2c1",
   885 => x"dbc27b75",
   886 => x"49bf97e8",
   887 => x"dcdbc21e",
   888 => x"d6d5c149",
   889 => x"7486c487",
   890 => x"ffc1c149",
   891 => x"c149c087",
   892 => x"c287dec3",
   893 => x"c048d0db",
   894 => x"dd49c178",
   895 => x"fd2687cb",
   896 => x"6f4c87ff",
   897 => x"6e696461",
   898 => x"2e2e2e67",
   899 => x"5b5e0e00",
   900 => x"4b710e5c",
   901 => x"d4dbc24a",
   902 => x"497282bf",
   903 => x"7087e6fc",
   904 => x"c4029c4c",
   905 => x"e9ec4987",
   906 => x"d4dbc287",
   907 => x"c178c048",
   908 => x"87d5dc49",
   909 => x"0e87ccfd",
   910 => x"5d5c5b5e",
   911 => x"c286f40e",
   912 => x"c04ddece",
   913 => x"48a6c44c",
   914 => x"dbc278c0",
   915 => x"c049bfd4",
   916 => x"c1c106a9",
   917 => x"decec287",
   918 => x"c0029848",
   919 => x"f2c087f8",
   920 => x"66c81ed7",
   921 => x"c487c702",
   922 => x"78c048a6",
   923 => x"a6c487c5",
   924 => x"c478c148",
   925 => x"d1ec4966",
   926 => x"7086c487",
   927 => x"c484c14d",
   928 => x"80c14866",
   929 => x"c258a6c8",
   930 => x"49bfd4db",
   931 => x"87c603ac",
   932 => x"ff059d75",
   933 => x"4cc087c8",
   934 => x"c3029d75",
   935 => x"f2c087e0",
   936 => x"66c81ed7",
   937 => x"cc87c702",
   938 => x"78c048a6",
   939 => x"a6cc87c5",
   940 => x"cc78c148",
   941 => x"d1eb4966",
   942 => x"7086c487",
   943 => x"c2026e7e",
   944 => x"496e87e9",
   945 => x"699781cb",
   946 => x"0299d049",
   947 => x"c087d6c1",
   948 => x"744acdf8",
   949 => x"c191cb49",
   950 => x"7281eed8",
   951 => x"c381c879",
   952 => x"497451ff",
   953 => x"dbc291de",
   954 => x"85714de9",
   955 => x"7d97c1c2",
   956 => x"c049a5c1",
   957 => x"d6c251e0",
   958 => x"02bf97ee",
   959 => x"84c187d2",
   960 => x"c24ba5c2",
   961 => x"db4aeed6",
   962 => x"dbc6ff49",
   963 => x"87dbc187",
   964 => x"c049a5cd",
   965 => x"c284c151",
   966 => x"4a6e4ba5",
   967 => x"c6ff49cb",
   968 => x"c6c187c6",
   969 => x"c9f6c087",
   970 => x"cb49744a",
   971 => x"eed8c191",
   972 => x"c2797281",
   973 => x"bf97eed6",
   974 => x"7487d802",
   975 => x"c191de49",
   976 => x"e9dbc284",
   977 => x"c283714b",
   978 => x"dd4aeed6",
   979 => x"d7c5ff49",
   980 => x"7487d887",
   981 => x"c293de4b",
   982 => x"cb83e9db",
   983 => x"51c049a3",
   984 => x"6e7384c1",
   985 => x"ff49cb4a",
   986 => x"c487fdc4",
   987 => x"80c14866",
   988 => x"c758a6c8",
   989 => x"c5c003ac",
   990 => x"fc056e87",
   991 => x"487487e0",
   992 => x"fcf78ef4",
   993 => x"1e731e87",
   994 => x"cb494b71",
   995 => x"eed8c191",
   996 => x"4aa1c881",
   997 => x"48cacdc2",
   998 => x"a1c95012",
   999 => x"c4f5c04a",
  1000 => x"ca501248",
  1001 => x"e8dbc281",
  1002 => x"c2501148",
  1003 => x"bf97e8db",
  1004 => x"49c01e49",
  1005 => x"87c3cec1",
  1006 => x"48d0dbc2",
  1007 => x"49c178de",
  1008 => x"2687c6d6",
  1009 => x"1e87fef6",
  1010 => x"cb494a71",
  1011 => x"eed8c191",
  1012 => x"1181c881",
  1013 => x"d4dbc248",
  1014 => x"d4dbc258",
  1015 => x"c178c048",
  1016 => x"87e5d549",
  1017 => x"c01e4f26",
  1018 => x"e4fbc049",
  1019 => x"1e4f2687",
  1020 => x"d2029971",
  1021 => x"c3dac187",
  1022 => x"f750c048",
  1023 => x"c7ffc080",
  1024 => x"e7d8c140",
  1025 => x"c187ce78",
  1026 => x"c148ffd9",
  1027 => x"fc78e0d8",
  1028 => x"e6ffc080",
  1029 => x"0e4f2678",
  1030 => x"0e5c5b5e",
  1031 => x"cb4a4c71",
  1032 => x"eed8c192",
  1033 => x"49a2c882",
  1034 => x"974ba2c9",
  1035 => x"971e4b6b",
  1036 => x"ca1e4969",
  1037 => x"c0491282",
  1038 => x"c087dfe6",
  1039 => x"87c9d449",
  1040 => x"f8c04974",
  1041 => x"8ef887e6",
  1042 => x"1e87f8f4",
  1043 => x"4b711e73",
  1044 => x"87c3ff49",
  1045 => x"fefe4973",
  1046 => x"87e9f487",
  1047 => x"711e731e",
  1048 => x"4aa3c64b",
  1049 => x"c187db02",
  1050 => x"87d6028a",
  1051 => x"dac1028a",
  1052 => x"c0028a87",
  1053 => x"028a87fc",
  1054 => x"8a87e1c0",
  1055 => x"c187cb02",
  1056 => x"49c787db",
  1057 => x"c187c0fd",
  1058 => x"dbc287de",
  1059 => x"c102bfd4",
  1060 => x"c14887cb",
  1061 => x"d8dbc288",
  1062 => x"87c1c158",
  1063 => x"bfd8dbc2",
  1064 => x"87f9c002",
  1065 => x"bfd4dbc2",
  1066 => x"c280c148",
  1067 => x"c058d8db",
  1068 => x"dbc287eb",
  1069 => x"c649bfd4",
  1070 => x"d8dbc289",
  1071 => x"a9b7c059",
  1072 => x"c287da03",
  1073 => x"c048d4db",
  1074 => x"c287d278",
  1075 => x"02bfd8db",
  1076 => x"dbc287cb",
  1077 => x"c648bfd4",
  1078 => x"d8dbc280",
  1079 => x"d149c058",
  1080 => x"497387e7",
  1081 => x"87c4f6c0",
  1082 => x"0e87daf2",
  1083 => x"0e5c5b5e",
  1084 => x"66cc4c71",
  1085 => x"cb4b741e",
  1086 => x"eed8c193",
  1087 => x"4aa3c483",
  1088 => x"fefe496a",
  1089 => x"fec087f2",
  1090 => x"a3c87bc5",
  1091 => x"5166d449",
  1092 => x"d849a3c9",
  1093 => x"a3ca5166",
  1094 => x"5166dc49",
  1095 => x"87e3f126",
  1096 => x"5c5b5e0e",
  1097 => x"d0ff0e5d",
  1098 => x"59a6d886",
  1099 => x"c048a6c4",
  1100 => x"c180c478",
  1101 => x"c47866c4",
  1102 => x"c478c180",
  1103 => x"c278c180",
  1104 => x"c148d8db",
  1105 => x"d0dbc278",
  1106 => x"a8de48bf",
  1107 => x"f387cb05",
  1108 => x"497087e5",
  1109 => x"ce59a6c8",
  1110 => x"ede887f8",
  1111 => x"87cfe987",
  1112 => x"7087dce8",
  1113 => x"acfbc04c",
  1114 => x"87d0c102",
  1115 => x"c10566d4",
  1116 => x"1ec087c2",
  1117 => x"c11ec11e",
  1118 => x"c01ee1da",
  1119 => x"87ebfd49",
  1120 => x"4a66d0c1",
  1121 => x"496a82c4",
  1122 => x"517481c7",
  1123 => x"1ed81ec1",
  1124 => x"81c8496a",
  1125 => x"d887ece8",
  1126 => x"66c4c186",
  1127 => x"01a8c048",
  1128 => x"a6c487c7",
  1129 => x"ce78c148",
  1130 => x"66c4c187",
  1131 => x"cc88c148",
  1132 => x"87c358a6",
  1133 => x"cc87f8e7",
  1134 => x"78c248a6",
  1135 => x"cd029c74",
  1136 => x"66c487cc",
  1137 => x"66c8c148",
  1138 => x"c1cd03a8",
  1139 => x"48a6d887",
  1140 => x"eae678c0",
  1141 => x"c14c7087",
  1142 => x"c205acd0",
  1143 => x"66d887d6",
  1144 => x"87cee97e",
  1145 => x"a6dc4970",
  1146 => x"87d3e659",
  1147 => x"ecc04c70",
  1148 => x"eac105ac",
  1149 => x"4966c487",
  1150 => x"c0c191cb",
  1151 => x"a1c48166",
  1152 => x"c84d6a4a",
  1153 => x"66d84aa1",
  1154 => x"c7ffc052",
  1155 => x"87efe579",
  1156 => x"029c4c70",
  1157 => x"fbc087d8",
  1158 => x"87d202ac",
  1159 => x"dee55574",
  1160 => x"9c4c7087",
  1161 => x"c087c702",
  1162 => x"ff05acfb",
  1163 => x"e0c087ee",
  1164 => x"55c1c255",
  1165 => x"d47d97c0",
  1166 => x"a96e4966",
  1167 => x"c487db05",
  1168 => x"66c84866",
  1169 => x"87ca04a8",
  1170 => x"c14866c4",
  1171 => x"58a6c880",
  1172 => x"66c887c8",
  1173 => x"cc88c148",
  1174 => x"e2e458a6",
  1175 => x"c14c7087",
  1176 => x"c805acd0",
  1177 => x"4866d087",
  1178 => x"a6d480c1",
  1179 => x"acd0c158",
  1180 => x"87eafd02",
  1181 => x"d448a6dc",
  1182 => x"66d87866",
  1183 => x"a866dc48",
  1184 => x"87dcc905",
  1185 => x"48a6e0c0",
  1186 => x"c478f0c0",
  1187 => x"7866cc80",
  1188 => x"78c080c4",
  1189 => x"c048747e",
  1190 => x"f0c088fb",
  1191 => x"987058a6",
  1192 => x"87d7c802",
  1193 => x"c088cb48",
  1194 => x"7058a6f0",
  1195 => x"e9c00298",
  1196 => x"88c94887",
  1197 => x"58a6f0c0",
  1198 => x"c3029870",
  1199 => x"c44887e1",
  1200 => x"a6f0c088",
  1201 => x"02987058",
  1202 => x"c14887d6",
  1203 => x"a6f0c088",
  1204 => x"02987058",
  1205 => x"c787c8c3",
  1206 => x"e0c087db",
  1207 => x"78c048a6",
  1208 => x"c14866cc",
  1209 => x"58a6d080",
  1210 => x"7087d4e2",
  1211 => x"acecc04c",
  1212 => x"c087d502",
  1213 => x"c60266e0",
  1214 => x"a6e4c087",
  1215 => x"7487c95c",
  1216 => x"88f0c048",
  1217 => x"58a6e8c0",
  1218 => x"02acecc0",
  1219 => x"eee187cc",
  1220 => x"c04c7087",
  1221 => x"ff05acec",
  1222 => x"e0c087f4",
  1223 => x"66d41e66",
  1224 => x"ecc01e49",
  1225 => x"dac11e66",
  1226 => x"66d41ee1",
  1227 => x"87fbf649",
  1228 => x"1eca1ec0",
  1229 => x"cb4966dc",
  1230 => x"66d8c191",
  1231 => x"48a6d881",
  1232 => x"d878a1c4",
  1233 => x"e149bf66",
  1234 => x"86d887f9",
  1235 => x"06a8b7c0",
  1236 => x"c187c7c1",
  1237 => x"c81ede1e",
  1238 => x"e149bf66",
  1239 => x"86c887e5",
  1240 => x"c0484970",
  1241 => x"e4c08808",
  1242 => x"b7c058a6",
  1243 => x"e9c006a8",
  1244 => x"66e0c087",
  1245 => x"a8b7dd48",
  1246 => x"6e87df03",
  1247 => x"e0c049bf",
  1248 => x"e0c08166",
  1249 => x"c1496651",
  1250 => x"81bf6e81",
  1251 => x"c051c1c2",
  1252 => x"c24966e0",
  1253 => x"81bf6e81",
  1254 => x"7ec151c0",
  1255 => x"e287dcc4",
  1256 => x"e4c087d0",
  1257 => x"c9e258a6",
  1258 => x"a6e8c087",
  1259 => x"a8ecc058",
  1260 => x"87cbc005",
  1261 => x"48a6e4c0",
  1262 => x"7866e0c0",
  1263 => x"ff87c4c0",
  1264 => x"c487fcde",
  1265 => x"91cb4966",
  1266 => x"4866c0c1",
  1267 => x"7e708071",
  1268 => x"82c84a6e",
  1269 => x"81ca496e",
  1270 => x"5166e0c0",
  1271 => x"4966e4c0",
  1272 => x"e0c081c1",
  1273 => x"48c18966",
  1274 => x"49703071",
  1275 => x"977189c1",
  1276 => x"c5dfc27a",
  1277 => x"e0c049bf",
  1278 => x"6a972966",
  1279 => x"9871484a",
  1280 => x"58a6f0c0",
  1281 => x"81c4496e",
  1282 => x"66dc4d69",
  1283 => x"a866d848",
  1284 => x"87c8c002",
  1285 => x"c048a6d8",
  1286 => x"87c5c078",
  1287 => x"c148a6d8",
  1288 => x"1e66d878",
  1289 => x"751ee0c0",
  1290 => x"d6deff49",
  1291 => x"7086c887",
  1292 => x"acb7c04c",
  1293 => x"87d4c106",
  1294 => x"e0c08574",
  1295 => x"75897449",
  1296 => x"c6d5c14b",
  1297 => x"f1fe714a",
  1298 => x"85c287de",
  1299 => x"4866e8c0",
  1300 => x"ecc080c1",
  1301 => x"ecc058a6",
  1302 => x"81c14966",
  1303 => x"c002a970",
  1304 => x"a6d887c8",
  1305 => x"c078c048",
  1306 => x"a6d887c5",
  1307 => x"d878c148",
  1308 => x"a4c21e66",
  1309 => x"48e0c049",
  1310 => x"49708871",
  1311 => x"ff49751e",
  1312 => x"c887c0dd",
  1313 => x"a8b7c086",
  1314 => x"87c0ff01",
  1315 => x"0266e8c0",
  1316 => x"6e87d1c0",
  1317 => x"c081c949",
  1318 => x"6e5166e8",
  1319 => x"d7c0c148",
  1320 => x"87ccc078",
  1321 => x"81c9496e",
  1322 => x"486e51c2",
  1323 => x"78cbc1c1",
  1324 => x"c6c07ec1",
  1325 => x"f6dbff87",
  1326 => x"6e4c7087",
  1327 => x"87f5c002",
  1328 => x"c84866c4",
  1329 => x"c004a866",
  1330 => x"66c487cb",
  1331 => x"c880c148",
  1332 => x"e0c058a6",
  1333 => x"4866c887",
  1334 => x"a6cc88c1",
  1335 => x"87d5c058",
  1336 => x"05acc6c1",
  1337 => x"cc87c8c0",
  1338 => x"80c14866",
  1339 => x"ff58a6d0",
  1340 => x"7087fcda",
  1341 => x"4866d04c",
  1342 => x"a6d480c1",
  1343 => x"029c7458",
  1344 => x"c487cbc0",
  1345 => x"c8c14866",
  1346 => x"f204a866",
  1347 => x"daff87ff",
  1348 => x"66c487d4",
  1349 => x"03a8c748",
  1350 => x"c287e5c0",
  1351 => x"c048d8db",
  1352 => x"4966c478",
  1353 => x"c0c191cb",
  1354 => x"a1c48166",
  1355 => x"c04a6a4a",
  1356 => x"66c47952",
  1357 => x"c880c148",
  1358 => x"a8c758a6",
  1359 => x"87dbff04",
  1360 => x"e08ed0ff",
  1361 => x"203a87fb",
  1362 => x"1e731e00",
  1363 => x"029b4b71",
  1364 => x"dbc287c6",
  1365 => x"78c048d4",
  1366 => x"dbc21ec7",
  1367 => x"1e49bfd4",
  1368 => x"1eeed8c1",
  1369 => x"bfd0dbc2",
  1370 => x"87f4ee49",
  1371 => x"dbc286cc",
  1372 => x"e949bfd0",
  1373 => x"9b7387f9",
  1374 => x"c187c802",
  1375 => x"c049eed8",
  1376 => x"ff87fbe4",
  1377 => x"1e87fedf",
  1378 => x"48cacdc2",
  1379 => x"dac150c0",
  1380 => x"c049bfd1",
  1381 => x"c087f7f2",
  1382 => x"1e4f2648",
  1383 => x"c187e1c7",
  1384 => x"87e5fe49",
  1385 => x"87fdf3fe",
  1386 => x"cd029870",
  1387 => x"d8fbfe87",
  1388 => x"02987087",
  1389 => x"4ac187c4",
  1390 => x"4ac087c2",
  1391 => x"ce059a72",
  1392 => x"c11ec087",
  1393 => x"c049ebd7",
  1394 => x"c487c1f0",
  1395 => x"c087fe86",
  1396 => x"f6d7c11e",
  1397 => x"f3efc049",
  1398 => x"fe1ec087",
  1399 => x"497087e9",
  1400 => x"87e8efc0",
  1401 => x"f887d8c3",
  1402 => x"534f268e",
  1403 => x"61662044",
  1404 => x"64656c69",
  1405 => x"6f42002e",
  1406 => x"6e69746f",
  1407 => x"2e2e2e67",
  1408 => x"e7c01e00",
  1409 => x"87fa87d4",
  1410 => x"c21e4f26",
  1411 => x"c048d4db",
  1412 => x"d0dbc278",
  1413 => x"fe78c048",
  1414 => x"87e587c1",
  1415 => x"4f2648c0",
  1416 => x"78452080",
  1417 => x"80007469",
  1418 => x"63614220",
  1419 => x"0fc7006b",
  1420 => x"26e90000",
  1421 => x"00000000",
  1422 => x"000fc700",
  1423 => x"00270700",
  1424 => x"00000000",
  1425 => x"00000fc7",
  1426 => x"00002725",
  1427 => x"c7000000",
  1428 => x"4300000f",
  1429 => x"00000027",
  1430 => x"0fc70000",
  1431 => x"27610000",
  1432 => x"00000000",
  1433 => x"000fc700",
  1434 => x"00277f00",
  1435 => x"00000000",
  1436 => x"00000fc7",
  1437 => x"0000279d",
  1438 => x"c7000000",
  1439 => x"0000000f",
  1440 => x"00000000",
  1441 => x"105c0000",
  1442 => x"00000000",
  1443 => x"00000000",
  1444 => x"00169500",
  1445 => x"4f4f4200",
  1446 => x"20202054",
  1447 => x"4d4f5220",
  1448 => x"616f4c00",
  1449 => x"2e2a2064",
  1450 => x"f0fe1e00",
  1451 => x"cd78c048",
  1452 => x"26097909",
  1453 => x"fe1e1e4f",
  1454 => x"487ebff0",
  1455 => x"1e4f2626",
  1456 => x"c148f0fe",
  1457 => x"1e4f2678",
  1458 => x"c048f0fe",
  1459 => x"1e4f2678",
  1460 => x"52c04a71",
  1461 => x"0e4f2652",
  1462 => x"5d5c5b5e",
  1463 => x"7186f40e",
  1464 => x"7e6d974d",
  1465 => x"974ca5c1",
  1466 => x"a6c8486c",
  1467 => x"c4486e58",
  1468 => x"c505a866",
  1469 => x"c048ff87",
  1470 => x"caff87e6",
  1471 => x"49a5c287",
  1472 => x"714b6c97",
  1473 => x"6b974ba3",
  1474 => x"7e6c974b",
  1475 => x"80c1486e",
  1476 => x"c758a6c8",
  1477 => x"58a6cc98",
  1478 => x"fe7c9770",
  1479 => x"487387e1",
  1480 => x"4d268ef4",
  1481 => x"4b264c26",
  1482 => x"5e0e4f26",
  1483 => x"f40e5c5b",
  1484 => x"d84c7186",
  1485 => x"ffc34a66",
  1486 => x"4ba4c29a",
  1487 => x"73496c97",
  1488 => x"517249a1",
  1489 => x"6e7e6c97",
  1490 => x"c880c148",
  1491 => x"98c758a6",
  1492 => x"7058a6cc",
  1493 => x"ff8ef454",
  1494 => x"1e1e87ca",
  1495 => x"e087e8fd",
  1496 => x"c0494abf",
  1497 => x"0299c0e0",
  1498 => x"1e7287cb",
  1499 => x"49fbdec2",
  1500 => x"c487f7fe",
  1501 => x"87fdfc86",
  1502 => x"c2fd7e70",
  1503 => x"4f262687",
  1504 => x"fbdec21e",
  1505 => x"87c7fd49",
  1506 => x"49daddc1",
  1507 => x"c487dafc",
  1508 => x"4f2687ff",
  1509 => x"5c5b5e0e",
  1510 => x"dfc20e5d",
  1511 => x"c14abfda",
  1512 => x"49bfe8df",
  1513 => x"71bc724c",
  1514 => x"87dbfc4d",
  1515 => x"49744bc0",
  1516 => x"d50299d0",
  1517 => x"d0497587",
  1518 => x"c01e7199",
  1519 => x"e0e5c11e",
  1520 => x"1282734a",
  1521 => x"87e4c049",
  1522 => x"2cc186c8",
  1523 => x"abc8832d",
  1524 => x"87daff04",
  1525 => x"c187e8fb",
  1526 => x"c248e8df",
  1527 => x"78bfdadf",
  1528 => x"4c264d26",
  1529 => x"4f264b26",
  1530 => x"00000000",
  1531 => x"48d0ff1e",
  1532 => x"ff78e1c8",
  1533 => x"78c548d4",
  1534 => x"c30266c4",
  1535 => x"78e0c387",
  1536 => x"c60266c8",
  1537 => x"48d4ff87",
  1538 => x"ff78f0c3",
  1539 => x"787148d4",
  1540 => x"c848d0ff",
  1541 => x"e0c078e1",
  1542 => x"1e4f2678",
  1543 => x"dec21e73",
  1544 => x"f2fa49fb",
  1545 => x"c04a7087",
  1546 => x"c204aab7",
  1547 => x"e0c387cd",
  1548 => x"87c905aa",
  1549 => x"48c4e3c1",
  1550 => x"fec178c1",
  1551 => x"aaf0c387",
  1552 => x"c187c905",
  1553 => x"c148c0e3",
  1554 => x"87dfc178",
  1555 => x"bfc4e3c1",
  1556 => x"7287c702",
  1557 => x"b3c0c24b",
  1558 => x"4b7287c2",
  1559 => x"bfc0e3c1",
  1560 => x"87e0c002",
  1561 => x"b7c44973",
  1562 => x"e4c19129",
  1563 => x"4a7381e0",
  1564 => x"92c29acf",
  1565 => x"307248c1",
  1566 => x"baff4a70",
  1567 => x"98694872",
  1568 => x"87db7970",
  1569 => x"b7c44973",
  1570 => x"e4c19129",
  1571 => x"4a7381e0",
  1572 => x"92c29acf",
  1573 => x"307248c3",
  1574 => x"69484a70",
  1575 => x"c17970b0",
  1576 => x"c048c4e3",
  1577 => x"c0e3c178",
  1578 => x"c278c048",
  1579 => x"f849fbde",
  1580 => x"4a7087e5",
  1581 => x"03aab7c0",
  1582 => x"c087f3fd",
  1583 => x"87e4fc48",
  1584 => x"00000000",
  1585 => x"00000000",
  1586 => x"494a711e",
  1587 => x"2687ccfd",
  1588 => x"4ac01e4f",
  1589 => x"91c44972",
  1590 => x"81e0e4c1",
  1591 => x"82c179c0",
  1592 => x"04aab7d0",
  1593 => x"4f2687ee",
  1594 => x"5c5b5e0e",
  1595 => x"4d710e5d",
  1596 => x"7587d4f7",
  1597 => x"2ab7c44a",
  1598 => x"e0e4c192",
  1599 => x"cf4c7582",
  1600 => x"6a94c29c",
  1601 => x"2b744b49",
  1602 => x"48c29bc3",
  1603 => x"4c703074",
  1604 => x"4874bcff",
  1605 => x"7a709871",
  1606 => x"7387e4f6",
  1607 => x"87c0fb48",
  1608 => x"00000000",
  1609 => x"00000000",
  1610 => x"00000000",
  1611 => x"00000000",
  1612 => x"00000000",
  1613 => x"00000000",
  1614 => x"00000000",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"00000000",
  1618 => x"00000000",
  1619 => x"00000000",
  1620 => x"00000000",
  1621 => x"00000000",
  1622 => x"00000000",
  1623 => x"00000000",
  1624 => x"25261e16",
  1625 => x"3e3d362e",
  1626 => x"48d0ff1e",
  1627 => x"7178e1c8",
  1628 => x"08d4ff48",
  1629 => x"4866c478",
  1630 => x"7808d4ff",
  1631 => x"711e4f26",
  1632 => x"4966c44a",
  1633 => x"ff49721e",
  1634 => x"d0ff87de",
  1635 => x"78e0c048",
  1636 => x"1e4f2626",
  1637 => x"b7c24a71",
  1638 => x"87c303aa",
  1639 => x"ce87c282",
  1640 => x"1e66c482",
  1641 => x"d5ff4972",
  1642 => x"4f262687",
  1643 => x"4ad4ff1e",
  1644 => x"ff7affc3",
  1645 => x"e1c848d0",
  1646 => x"c27ade78",
  1647 => x"7abfc5df",
  1648 => x"28c84849",
  1649 => x"48717a70",
  1650 => x"7a7028d0",
  1651 => x"28d84871",
  1652 => x"d0ff7a70",
  1653 => x"78e0c048",
  1654 => x"5e0e4f26",
  1655 => x"0e5d5c5b",
  1656 => x"dfc24c71",
  1657 => x"4b4dbfc5",
  1658 => x"66d02b74",
  1659 => x"d483c19b",
  1660 => x"c204ab66",
  1661 => x"744bc087",
  1662 => x"4966d04a",
  1663 => x"b9ff3172",
  1664 => x"48739975",
  1665 => x"4a703072",
  1666 => x"c2b07148",
  1667 => x"fe58c9df",
  1668 => x"4d2687da",
  1669 => x"4b264c26",
  1670 => x"ff1e4f26",
  1671 => x"c9c848d0",
  1672 => x"ff487178",
  1673 => x"267808d4",
  1674 => x"4a711e4f",
  1675 => x"ff87eb49",
  1676 => x"78c848d0",
  1677 => x"731e4f26",
  1678 => x"c24b711e",
  1679 => x"02bfd5df",
  1680 => x"ebc287c3",
  1681 => x"48d0ff87",
  1682 => x"7378c9c8",
  1683 => x"b1e0c049",
  1684 => x"7148d4ff",
  1685 => x"c9dfc278",
  1686 => x"c878c048",
  1687 => x"87c50266",
  1688 => x"c249ffc3",
  1689 => x"c249c087",
  1690 => x"cc59d1df",
  1691 => x"87c60266",
  1692 => x"4ad5d5c5",
  1693 => x"ffcf87c4",
  1694 => x"dfc24aff",
  1695 => x"dfc25ad5",
  1696 => x"78c148d5",
  1697 => x"4d2687c4",
  1698 => x"4b264c26",
  1699 => x"5e0e4f26",
  1700 => x"0e5d5c5b",
  1701 => x"dfc24a71",
  1702 => x"724cbfd1",
  1703 => x"87cb029a",
  1704 => x"c191c849",
  1705 => x"714bece8",
  1706 => x"c187c483",
  1707 => x"c04becec",
  1708 => x"7449134d",
  1709 => x"cddfc299",
  1710 => x"d4ffb9bf",
  1711 => x"c1787148",
  1712 => x"c8852cb7",
  1713 => x"e804adb7",
  1714 => x"c9dfc287",
  1715 => x"80c848bf",
  1716 => x"58cddfc2",
  1717 => x"1e87effe",
  1718 => x"4b711e73",
  1719 => x"029a4a13",
  1720 => x"497287cb",
  1721 => x"1387e7fe",
  1722 => x"f5059a4a",
  1723 => x"87dafe87",
  1724 => x"c9dfc21e",
  1725 => x"dfc249bf",
  1726 => x"a1c148c9",
  1727 => x"b7c0c478",
  1728 => x"87db03a9",
  1729 => x"c248d4ff",
  1730 => x"78bfcddf",
  1731 => x"bfc9dfc2",
  1732 => x"c9dfc249",
  1733 => x"78a1c148",
  1734 => x"a9b7c0c4",
  1735 => x"ff87e504",
  1736 => x"78c848d0",
  1737 => x"48d5dfc2",
  1738 => x"4f2678c0",
  1739 => x"00000000",
  1740 => x"00000000",
  1741 => x"5f000000",
  1742 => x"0000005f",
  1743 => x"00030300",
  1744 => x"00000303",
  1745 => x"147f7f14",
  1746 => x"00147f7f",
  1747 => x"6b2e2400",
  1748 => x"00123a6b",
  1749 => x"18366a4c",
  1750 => x"0032566c",
  1751 => x"594f7e30",
  1752 => x"40683a77",
  1753 => x"07040000",
  1754 => x"00000003",
  1755 => x"3e1c0000",
  1756 => x"00004163",
  1757 => x"63410000",
  1758 => x"00001c3e",
  1759 => x"1c3e2a08",
  1760 => x"082a3e1c",
  1761 => x"3e080800",
  1762 => x"0008083e",
  1763 => x"e0800000",
  1764 => x"00000060",
  1765 => x"08080800",
  1766 => x"00080808",
  1767 => x"60000000",
  1768 => x"00000060",
  1769 => x"18306040",
  1770 => x"0103060c",
  1771 => x"597f3e00",
  1772 => x"003e7f4d",
  1773 => x"7f060400",
  1774 => x"0000007f",
  1775 => x"71634200",
  1776 => x"00464f59",
  1777 => x"49632200",
  1778 => x"00367f49",
  1779 => x"13161c18",
  1780 => x"00107f7f",
  1781 => x"45672700",
  1782 => x"00397d45",
  1783 => x"4b7e3c00",
  1784 => x"00307949",
  1785 => x"71010100",
  1786 => x"00070f79",
  1787 => x"497f3600",
  1788 => x"00367f49",
  1789 => x"494f0600",
  1790 => x"001e3f69",
  1791 => x"66000000",
  1792 => x"00000066",
  1793 => x"e6800000",
  1794 => x"00000066",
  1795 => x"14080800",
  1796 => x"00222214",
  1797 => x"14141400",
  1798 => x"00141414",
  1799 => x"14222200",
  1800 => x"00080814",
  1801 => x"51030200",
  1802 => x"00060f59",
  1803 => x"5d417f3e",
  1804 => x"001e1f55",
  1805 => x"097f7e00",
  1806 => x"007e7f09",
  1807 => x"497f7f00",
  1808 => x"00367f49",
  1809 => x"633e1c00",
  1810 => x"00414141",
  1811 => x"417f7f00",
  1812 => x"001c3e63",
  1813 => x"497f7f00",
  1814 => x"00414149",
  1815 => x"097f7f00",
  1816 => x"00010109",
  1817 => x"417f3e00",
  1818 => x"007a7b49",
  1819 => x"087f7f00",
  1820 => x"007f7f08",
  1821 => x"7f410000",
  1822 => x"0000417f",
  1823 => x"40602000",
  1824 => x"003f7f40",
  1825 => x"1c087f7f",
  1826 => x"00416336",
  1827 => x"407f7f00",
  1828 => x"00404040",
  1829 => x"0c067f7f",
  1830 => x"007f7f06",
  1831 => x"0c067f7f",
  1832 => x"007f7f18",
  1833 => x"417f3e00",
  1834 => x"003e7f41",
  1835 => x"097f7f00",
  1836 => x"00060f09",
  1837 => x"61417f3e",
  1838 => x"00407e7f",
  1839 => x"097f7f00",
  1840 => x"00667f19",
  1841 => x"4d6f2600",
  1842 => x"00327b59",
  1843 => x"7f010100",
  1844 => x"0001017f",
  1845 => x"407f3f00",
  1846 => x"003f7f40",
  1847 => x"703f0f00",
  1848 => x"000f3f70",
  1849 => x"18307f7f",
  1850 => x"007f7f30",
  1851 => x"1c366341",
  1852 => x"4163361c",
  1853 => x"7c060301",
  1854 => x"0103067c",
  1855 => x"4d597161",
  1856 => x"00414347",
  1857 => x"7f7f0000",
  1858 => x"00004141",
  1859 => x"0c060301",
  1860 => x"40603018",
  1861 => x"41410000",
  1862 => x"00007f7f",
  1863 => x"03060c08",
  1864 => x"00080c06",
  1865 => x"80808080",
  1866 => x"00808080",
  1867 => x"03000000",
  1868 => x"00000407",
  1869 => x"54742000",
  1870 => x"00787c54",
  1871 => x"447f7f00",
  1872 => x"00387c44",
  1873 => x"447c3800",
  1874 => x"00004444",
  1875 => x"447c3800",
  1876 => x"007f7f44",
  1877 => x"547c3800",
  1878 => x"00185c54",
  1879 => x"7f7e0400",
  1880 => x"00000505",
  1881 => x"a4bc1800",
  1882 => x"007cfca4",
  1883 => x"047f7f00",
  1884 => x"00787c04",
  1885 => x"3d000000",
  1886 => x"0000407d",
  1887 => x"80808000",
  1888 => x"00007dfd",
  1889 => x"107f7f00",
  1890 => x"00446c38",
  1891 => x"3f000000",
  1892 => x"0000407f",
  1893 => x"180c7c7c",
  1894 => x"00787c0c",
  1895 => x"047c7c00",
  1896 => x"00787c04",
  1897 => x"447c3800",
  1898 => x"00387c44",
  1899 => x"24fcfc00",
  1900 => x"00183c24",
  1901 => x"243c1800",
  1902 => x"00fcfc24",
  1903 => x"047c7c00",
  1904 => x"00080c04",
  1905 => x"545c4800",
  1906 => x"00207454",
  1907 => x"7f3f0400",
  1908 => x"00004444",
  1909 => x"407c3c00",
  1910 => x"007c7c40",
  1911 => x"603c1c00",
  1912 => x"001c3c60",
  1913 => x"30607c3c",
  1914 => x"003c7c60",
  1915 => x"10386c44",
  1916 => x"00446c38",
  1917 => x"e0bc1c00",
  1918 => x"001c3c60",
  1919 => x"74644400",
  1920 => x"00444c5c",
  1921 => x"3e080800",
  1922 => x"00414177",
  1923 => x"7f000000",
  1924 => x"0000007f",
  1925 => x"77414100",
  1926 => x"0008083e",
  1927 => x"03010102",
  1928 => x"00010202",
  1929 => x"7f7f7f7f",
  1930 => x"007f7f7f",
  1931 => x"1c1c0808",
  1932 => x"7f7f3e3e",
  1933 => x"3e3e7f7f",
  1934 => x"08081c1c",
  1935 => x"7c181000",
  1936 => x"0010187c",
  1937 => x"7c301000",
  1938 => x"0010307c",
  1939 => x"60603010",
  1940 => x"00061e78",
  1941 => x"183c6642",
  1942 => x"0042663c",
  1943 => x"c26a3878",
  1944 => x"00386cc6",
  1945 => x"60000060",
  1946 => x"00600000",
  1947 => x"5c5b5e0e",
  1948 => x"711e0e5d",
  1949 => x"e6dfc24c",
  1950 => x"4bc04dbf",
  1951 => x"ab741ec0",
  1952 => x"c487c702",
  1953 => x"78c048a6",
  1954 => x"a6c487c5",
  1955 => x"c478c148",
  1956 => x"49731e66",
  1957 => x"c887dfee",
  1958 => x"49e0c086",
  1959 => x"c487efef",
  1960 => x"496a4aa5",
  1961 => x"f187f0f0",
  1962 => x"85cb87c6",
  1963 => x"b7c883c1",
  1964 => x"c7ff04ab",
  1965 => x"4d262687",
  1966 => x"4b264c26",
  1967 => x"711e4f26",
  1968 => x"eadfc24a",
  1969 => x"eadfc25a",
  1970 => x"4978c748",
  1971 => x"2687ddfe",
  1972 => x"1e731e4f",
  1973 => x"b7c04a71",
  1974 => x"87d303aa",
  1975 => x"bfe1c8c2",
  1976 => x"c187c405",
  1977 => x"c087c24b",
  1978 => x"e5c8c24b",
  1979 => x"c287c45b",
  1980 => x"c25ae5c8",
  1981 => x"4abfe1c8",
  1982 => x"c0c19ac1",
  1983 => x"e8ec49a2",
  1984 => x"c248fc87",
  1985 => x"78bfe1c8",
  1986 => x"1e87effe",
  1987 => x"66c44a71",
  1988 => x"e949721e",
  1989 => x"262687fd",
  1990 => x"c8c21e4f",
  1991 => x"e649bfe1",
  1992 => x"dfc287e6",
  1993 => x"bfe848de",
  1994 => x"dadfc278",
  1995 => x"78bfec48",
  1996 => x"bfdedfc2",
  1997 => x"ffc3494a",
  1998 => x"2ab7c899",
  1999 => x"b0714872",
  2000 => x"58e6dfc2",
  2001 => x"5e0e4f26",
  2002 => x"0e5d5c5b",
  2003 => x"c8ff4b71",
  2004 => x"d9dfc287",
  2005 => x"7350c048",
  2006 => x"87cce649",
  2007 => x"c24c4970",
  2008 => x"49eecb9c",
  2009 => x"7087c2cb",
  2010 => x"dfc24d49",
  2011 => x"05bf97d9",
  2012 => x"d087e2c1",
  2013 => x"dfc24966",
  2014 => x"0599bfe2",
  2015 => x"66d487d6",
  2016 => x"dadfc249",
  2017 => x"cb0599bf",
  2018 => x"e5497387",
  2019 => x"987087da",
  2020 => x"87c1c102",
  2021 => x"c0fe4cc1",
  2022 => x"ca497587",
  2023 => x"987087d7",
  2024 => x"c287c602",
  2025 => x"c148d9df",
  2026 => x"d9dfc250",
  2027 => x"c005bf97",
  2028 => x"dfc287e3",
  2029 => x"d049bfe2",
  2030 => x"ff059966",
  2031 => x"dfc287d6",
  2032 => x"d449bfda",
  2033 => x"ff059966",
  2034 => x"497387ca",
  2035 => x"7087d9e4",
  2036 => x"fffe0598",
  2037 => x"fb487487",
  2038 => x"5e0e87dc",
  2039 => x"0e5d5c5b",
  2040 => x"4dc086f4",
  2041 => x"7ebfec4c",
  2042 => x"c248a6c4",
  2043 => x"78bfe6df",
  2044 => x"1ec01ec1",
  2045 => x"cdfd49c7",
  2046 => x"7086c887",
  2047 => x"87cd0298",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
