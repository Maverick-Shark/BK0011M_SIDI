
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"e0",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"c4",x"e0",x"c2"),
    14 => (x"48",x"f8",x"cd",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ff",x"d6"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"d4",x"ff",x"1e",x"4f"),
    50 => (x"78",x"ff",x"c3",x"48"),
    51 => (x"66",x"c4",x"51",x"68"),
    52 => (x"c8",x"88",x"c1",x"48"),
    53 => (x"98",x"70",x"58",x"a6"),
    54 => (x"26",x"87",x"eb",x"05"),
    55 => (x"1e",x"73",x"1e",x"4f"),
    56 => (x"c3",x"4b",x"d4",x"ff"),
    57 => (x"4a",x"6b",x"7b",x"ff"),
    58 => (x"6b",x"7b",x"ff",x"c3"),
    59 => (x"72",x"32",x"c8",x"49"),
    60 => (x"7b",x"ff",x"c3",x"b1"),
    61 => (x"31",x"c8",x"4a",x"6b"),
    62 => (x"ff",x"c3",x"b2",x"71"),
    63 => (x"c8",x"49",x"6b",x"7b"),
    64 => (x"71",x"b1",x"72",x"32"),
    65 => (x"26",x"87",x"c4",x"48"),
    66 => (x"26",x"4c",x"26",x"4d"),
    67 => (x"0e",x"4f",x"26",x"4b"),
    68 => (x"5d",x"5c",x"5b",x"5e"),
    69 => (x"ff",x"4a",x"71",x"0e"),
    70 => (x"49",x"72",x"4c",x"d4"),
    71 => (x"71",x"99",x"ff",x"c3"),
    72 => (x"f8",x"cd",x"c2",x"7c"),
    73 => (x"87",x"c8",x"05",x"bf"),
    74 => (x"c9",x"48",x"66",x"d0"),
    75 => (x"58",x"a6",x"d4",x"30"),
    76 => (x"d8",x"49",x"66",x"d0"),
    77 => (x"99",x"ff",x"c3",x"29"),
    78 => (x"66",x"d0",x"7c",x"71"),
    79 => (x"c3",x"29",x"d0",x"49"),
    80 => (x"7c",x"71",x"99",x"ff"),
    81 => (x"c8",x"49",x"66",x"d0"),
    82 => (x"99",x"ff",x"c3",x"29"),
    83 => (x"66",x"d0",x"7c",x"71"),
    84 => (x"99",x"ff",x"c3",x"49"),
    85 => (x"49",x"72",x"7c",x"71"),
    86 => (x"ff",x"c3",x"29",x"d0"),
    87 => (x"6c",x"7c",x"71",x"99"),
    88 => (x"ff",x"f0",x"c9",x"4b"),
    89 => (x"ab",x"ff",x"c3",x"4d"),
    90 => (x"c3",x"87",x"d0",x"05"),
    91 => (x"4b",x"6c",x"7c",x"ff"),
    92 => (x"c6",x"02",x"8d",x"c1"),
    93 => (x"ab",x"ff",x"c3",x"87"),
    94 => (x"73",x"87",x"f0",x"02"),
    95 => (x"87",x"c7",x"fe",x"48"),
    96 => (x"ff",x"49",x"c0",x"1e"),
    97 => (x"ff",x"c3",x"48",x"d4"),
    98 => (x"c3",x"81",x"c1",x"78"),
    99 => (x"04",x"a9",x"b7",x"c8"),
   100 => (x"4f",x"26",x"87",x"f1"),
   101 => (x"e7",x"1e",x"73",x"1e"),
   102 => (x"df",x"f8",x"c4",x"87"),
   103 => (x"c0",x"1e",x"c0",x"4b"),
   104 => (x"f7",x"c1",x"f0",x"ff"),
   105 => (x"87",x"e7",x"fd",x"49"),
   106 => (x"a8",x"c1",x"86",x"c4"),
   107 => (x"87",x"ea",x"c0",x"05"),
   108 => (x"c3",x"48",x"d4",x"ff"),
   109 => (x"c0",x"c1",x"78",x"ff"),
   110 => (x"c0",x"c0",x"c0",x"c0"),
   111 => (x"f0",x"e1",x"c0",x"1e"),
   112 => (x"fd",x"49",x"e9",x"c1"),
   113 => (x"86",x"c4",x"87",x"c9"),
   114 => (x"ca",x"05",x"98",x"70"),
   115 => (x"48",x"d4",x"ff",x"87"),
   116 => (x"c1",x"78",x"ff",x"c3"),
   117 => (x"fe",x"87",x"cb",x"48"),
   118 => (x"8b",x"c1",x"87",x"e6"),
   119 => (x"87",x"fd",x"fe",x"05"),
   120 => (x"e6",x"fc",x"48",x"c0"),
   121 => (x"1e",x"73",x"1e",x"87"),
   122 => (x"c3",x"48",x"d4",x"ff"),
   123 => (x"4b",x"d3",x"78",x"ff"),
   124 => (x"ff",x"c0",x"1e",x"c0"),
   125 => (x"49",x"c1",x"c1",x"f0"),
   126 => (x"c4",x"87",x"d4",x"fc"),
   127 => (x"05",x"98",x"70",x"86"),
   128 => (x"d4",x"ff",x"87",x"ca"),
   129 => (x"78",x"ff",x"c3",x"48"),
   130 => (x"87",x"cb",x"48",x"c1"),
   131 => (x"c1",x"87",x"f1",x"fd"),
   132 => (x"db",x"ff",x"05",x"8b"),
   133 => (x"fb",x"48",x"c0",x"87"),
   134 => (x"5e",x"0e",x"87",x"f1"),
   135 => (x"ff",x"0e",x"5c",x"5b"),
   136 => (x"db",x"fd",x"4c",x"d4"),
   137 => (x"1e",x"ea",x"c6",x"87"),
   138 => (x"c1",x"f0",x"e1",x"c0"),
   139 => (x"de",x"fb",x"49",x"c8"),
   140 => (x"c1",x"86",x"c4",x"87"),
   141 => (x"87",x"c8",x"02",x"a8"),
   142 => (x"c0",x"87",x"ea",x"fe"),
   143 => (x"87",x"e2",x"c1",x"48"),
   144 => (x"70",x"87",x"da",x"fa"),
   145 => (x"ff",x"ff",x"cf",x"49"),
   146 => (x"a9",x"ea",x"c6",x"99"),
   147 => (x"fe",x"87",x"c8",x"02"),
   148 => (x"48",x"c0",x"87",x"d3"),
   149 => (x"c3",x"87",x"cb",x"c1"),
   150 => (x"f1",x"c0",x"7c",x"ff"),
   151 => (x"87",x"f4",x"fc",x"4b"),
   152 => (x"c0",x"02",x"98",x"70"),
   153 => (x"1e",x"c0",x"87",x"eb"),
   154 => (x"c1",x"f0",x"ff",x"c0"),
   155 => (x"de",x"fa",x"49",x"fa"),
   156 => (x"70",x"86",x"c4",x"87"),
   157 => (x"87",x"d9",x"05",x"98"),
   158 => (x"6c",x"7c",x"ff",x"c3"),
   159 => (x"7c",x"ff",x"c3",x"49"),
   160 => (x"c1",x"7c",x"7c",x"7c"),
   161 => (x"c4",x"02",x"99",x"c0"),
   162 => (x"d5",x"48",x"c1",x"87"),
   163 => (x"d1",x"48",x"c0",x"87"),
   164 => (x"05",x"ab",x"c2",x"87"),
   165 => (x"48",x"c0",x"87",x"c4"),
   166 => (x"8b",x"c1",x"87",x"c8"),
   167 => (x"87",x"fd",x"fe",x"05"),
   168 => (x"e4",x"f9",x"48",x"c0"),
   169 => (x"1e",x"73",x"1e",x"87"),
   170 => (x"48",x"f8",x"cd",x"c2"),
   171 => (x"4b",x"c7",x"78",x"c1"),
   172 => (x"c2",x"48",x"d0",x"ff"),
   173 => (x"87",x"c8",x"fb",x"78"),
   174 => (x"c3",x"48",x"d0",x"ff"),
   175 => (x"c0",x"1e",x"c0",x"78"),
   176 => (x"c0",x"c1",x"d0",x"e5"),
   177 => (x"87",x"c7",x"f9",x"49"),
   178 => (x"a8",x"c1",x"86",x"c4"),
   179 => (x"4b",x"87",x"c1",x"05"),
   180 => (x"c5",x"05",x"ab",x"c2"),
   181 => (x"c0",x"48",x"c0",x"87"),
   182 => (x"8b",x"c1",x"87",x"f9"),
   183 => (x"87",x"d0",x"ff",x"05"),
   184 => (x"c2",x"87",x"f7",x"fc"),
   185 => (x"70",x"58",x"fc",x"cd"),
   186 => (x"87",x"cd",x"05",x"98"),
   187 => (x"ff",x"c0",x"1e",x"c1"),
   188 => (x"49",x"d0",x"c1",x"f0"),
   189 => (x"c4",x"87",x"d8",x"f8"),
   190 => (x"48",x"d4",x"ff",x"86"),
   191 => (x"c2",x"78",x"ff",x"c3"),
   192 => (x"ce",x"c2",x"87",x"fe"),
   193 => (x"d0",x"ff",x"58",x"c0"),
   194 => (x"ff",x"78",x"c2",x"48"),
   195 => (x"ff",x"c3",x"48",x"d4"),
   196 => (x"f7",x"48",x"c1",x"78"),
   197 => (x"ff",x"1e",x"87",x"f5"),
   198 => (x"d0",x"ff",x"4a",x"d4"),
   199 => (x"78",x"d1",x"c4",x"48"),
   200 => (x"c1",x"7a",x"ff",x"c3"),
   201 => (x"87",x"f8",x"05",x"89"),
   202 => (x"73",x"1e",x"4f",x"26"),
   203 => (x"c5",x"4b",x"71",x"1e"),
   204 => (x"4a",x"df",x"cd",x"ee"),
   205 => (x"c3",x"48",x"d4",x"ff"),
   206 => (x"48",x"68",x"78",x"ff"),
   207 => (x"02",x"a8",x"fe",x"c3"),
   208 => (x"8a",x"c1",x"87",x"c5"),
   209 => (x"72",x"87",x"ed",x"05"),
   210 => (x"87",x"c5",x"05",x"9a"),
   211 => (x"ea",x"c0",x"48",x"c0"),
   212 => (x"02",x"9b",x"73",x"87"),
   213 => (x"66",x"c8",x"87",x"cc"),
   214 => (x"f5",x"49",x"73",x"1e"),
   215 => (x"86",x"c4",x"87",x"e7"),
   216 => (x"66",x"c8",x"87",x"c6"),
   217 => (x"87",x"ee",x"fe",x"49"),
   218 => (x"c3",x"48",x"d4",x"ff"),
   219 => (x"73",x"78",x"78",x"ff"),
   220 => (x"87",x"c5",x"05",x"9b"),
   221 => (x"d0",x"48",x"d0",x"ff"),
   222 => (x"f6",x"48",x"c1",x"78"),
   223 => (x"73",x"1e",x"87",x"cd"),
   224 => (x"c0",x"4a",x"71",x"1e"),
   225 => (x"48",x"d4",x"ff",x"4b"),
   226 => (x"ff",x"78",x"ff",x"c3"),
   227 => (x"c3",x"c4",x"48",x"d0"),
   228 => (x"48",x"d4",x"ff",x"78"),
   229 => (x"72",x"78",x"ff",x"c3"),
   230 => (x"f0",x"ff",x"c0",x"1e"),
   231 => (x"f5",x"49",x"d1",x"c1"),
   232 => (x"86",x"c4",x"87",x"ed"),
   233 => (x"cd",x"05",x"98",x"70"),
   234 => (x"1e",x"c0",x"c8",x"87"),
   235 => (x"fd",x"49",x"66",x"cc"),
   236 => (x"86",x"c4",x"87",x"f8"),
   237 => (x"d0",x"ff",x"4b",x"70"),
   238 => (x"73",x"78",x"c2",x"48"),
   239 => (x"87",x"cb",x"f5",x"48"),
   240 => (x"5c",x"5b",x"5e",x"0e"),
   241 => (x"1e",x"c0",x"0e",x"5d"),
   242 => (x"c1",x"f0",x"ff",x"c0"),
   243 => (x"fe",x"f4",x"49",x"c9"),
   244 => (x"c2",x"1e",x"d2",x"87"),
   245 => (x"fd",x"49",x"c0",x"ce"),
   246 => (x"86",x"c8",x"87",x"d0"),
   247 => (x"84",x"c1",x"4c",x"c0"),
   248 => (x"04",x"ac",x"b7",x"d2"),
   249 => (x"ce",x"c2",x"87",x"f8"),
   250 => (x"49",x"bf",x"97",x"c0"),
   251 => (x"c1",x"99",x"c0",x"c3"),
   252 => (x"c0",x"05",x"a9",x"c0"),
   253 => (x"ce",x"c2",x"87",x"e7"),
   254 => (x"49",x"bf",x"97",x"c7"),
   255 => (x"ce",x"c2",x"31",x"d0"),
   256 => (x"4a",x"bf",x"97",x"c8"),
   257 => (x"b1",x"72",x"32",x"c8"),
   258 => (x"97",x"c9",x"ce",x"c2"),
   259 => (x"71",x"b1",x"4a",x"bf"),
   260 => (x"ff",x"ff",x"cf",x"4c"),
   261 => (x"84",x"c1",x"9c",x"ff"),
   262 => (x"e7",x"c1",x"34",x"ca"),
   263 => (x"c9",x"ce",x"c2",x"87"),
   264 => (x"c1",x"49",x"bf",x"97"),
   265 => (x"c2",x"99",x"c6",x"31"),
   266 => (x"bf",x"97",x"ca",x"ce"),
   267 => (x"2a",x"b7",x"c7",x"4a"),
   268 => (x"ce",x"c2",x"b1",x"72"),
   269 => (x"4a",x"bf",x"97",x"c5"),
   270 => (x"c2",x"9d",x"cf",x"4d"),
   271 => (x"bf",x"97",x"c6",x"ce"),
   272 => (x"ca",x"9a",x"c3",x"4a"),
   273 => (x"c7",x"ce",x"c2",x"32"),
   274 => (x"c2",x"4b",x"bf",x"97"),
   275 => (x"c2",x"b2",x"73",x"33"),
   276 => (x"bf",x"97",x"c8",x"ce"),
   277 => (x"9b",x"c0",x"c3",x"4b"),
   278 => (x"73",x"2b",x"b7",x"c6"),
   279 => (x"c1",x"81",x"c2",x"b2"),
   280 => (x"70",x"30",x"71",x"48"),
   281 => (x"75",x"48",x"c1",x"49"),
   282 => (x"72",x"4d",x"70",x"30"),
   283 => (x"71",x"84",x"c1",x"4c"),
   284 => (x"b7",x"c0",x"c8",x"94"),
   285 => (x"87",x"cc",x"06",x"ad"),
   286 => (x"2d",x"b7",x"34",x"c1"),
   287 => (x"ad",x"b7",x"c0",x"c8"),
   288 => (x"87",x"f4",x"ff",x"01"),
   289 => (x"fe",x"f1",x"48",x"74"),
   290 => (x"5b",x"5e",x"0e",x"87"),
   291 => (x"f8",x"0e",x"5d",x"5c"),
   292 => (x"e6",x"d6",x"c2",x"86"),
   293 => (x"c2",x"78",x"c0",x"48"),
   294 => (x"c0",x"1e",x"de",x"ce"),
   295 => (x"87",x"de",x"fb",x"49"),
   296 => (x"98",x"70",x"86",x"c4"),
   297 => (x"c0",x"87",x"c5",x"05"),
   298 => (x"87",x"ce",x"c9",x"48"),
   299 => (x"7e",x"c1",x"4d",x"c0"),
   300 => (x"bf",x"e9",x"ed",x"c0"),
   301 => (x"d4",x"cf",x"c2",x"49"),
   302 => (x"4b",x"c8",x"71",x"4a"),
   303 => (x"70",x"87",x"eb",x"ee"),
   304 => (x"87",x"c2",x"05",x"98"),
   305 => (x"ed",x"c0",x"7e",x"c0"),
   306 => (x"c2",x"49",x"bf",x"e5"),
   307 => (x"71",x"4a",x"f0",x"cf"),
   308 => (x"d5",x"ee",x"4b",x"c8"),
   309 => (x"05",x"98",x"70",x"87"),
   310 => (x"7e",x"c0",x"87",x"c2"),
   311 => (x"fd",x"c0",x"02",x"6e"),
   312 => (x"e4",x"d5",x"c2",x"87"),
   313 => (x"d6",x"c2",x"4d",x"bf"),
   314 => (x"7e",x"bf",x"9f",x"dc"),
   315 => (x"ea",x"d6",x"c5",x"48"),
   316 => (x"87",x"c7",x"05",x"a8"),
   317 => (x"bf",x"e4",x"d5",x"c2"),
   318 => (x"6e",x"87",x"ce",x"4d"),
   319 => (x"d5",x"e9",x"ca",x"48"),
   320 => (x"87",x"c5",x"02",x"a8"),
   321 => (x"f1",x"c7",x"48",x"c0"),
   322 => (x"de",x"ce",x"c2",x"87"),
   323 => (x"f9",x"49",x"75",x"1e"),
   324 => (x"86",x"c4",x"87",x"ec"),
   325 => (x"c5",x"05",x"98",x"70"),
   326 => (x"c7",x"48",x"c0",x"87"),
   327 => (x"ed",x"c0",x"87",x"dc"),
   328 => (x"c2",x"49",x"bf",x"e5"),
   329 => (x"71",x"4a",x"f0",x"cf"),
   330 => (x"fd",x"ec",x"4b",x"c8"),
   331 => (x"05",x"98",x"70",x"87"),
   332 => (x"d6",x"c2",x"87",x"c8"),
   333 => (x"78",x"c1",x"48",x"e6"),
   334 => (x"ed",x"c0",x"87",x"da"),
   335 => (x"c2",x"49",x"bf",x"e9"),
   336 => (x"71",x"4a",x"d4",x"cf"),
   337 => (x"e1",x"ec",x"4b",x"c8"),
   338 => (x"02",x"98",x"70",x"87"),
   339 => (x"c0",x"87",x"c5",x"c0"),
   340 => (x"87",x"e6",x"c6",x"48"),
   341 => (x"97",x"dc",x"d6",x"c2"),
   342 => (x"d5",x"c1",x"49",x"bf"),
   343 => (x"cd",x"c0",x"05",x"a9"),
   344 => (x"dd",x"d6",x"c2",x"87"),
   345 => (x"c2",x"49",x"bf",x"97"),
   346 => (x"c0",x"02",x"a9",x"ea"),
   347 => (x"48",x"c0",x"87",x"c5"),
   348 => (x"c2",x"87",x"c7",x"c6"),
   349 => (x"bf",x"97",x"de",x"ce"),
   350 => (x"e9",x"c3",x"48",x"7e"),
   351 => (x"ce",x"c0",x"02",x"a8"),
   352 => (x"c3",x"48",x"6e",x"87"),
   353 => (x"c0",x"02",x"a8",x"eb"),
   354 => (x"48",x"c0",x"87",x"c5"),
   355 => (x"c2",x"87",x"eb",x"c5"),
   356 => (x"bf",x"97",x"e9",x"ce"),
   357 => (x"c0",x"05",x"99",x"49"),
   358 => (x"ce",x"c2",x"87",x"cc"),
   359 => (x"49",x"bf",x"97",x"ea"),
   360 => (x"c0",x"02",x"a9",x"c2"),
   361 => (x"48",x"c0",x"87",x"c5"),
   362 => (x"c2",x"87",x"cf",x"c5"),
   363 => (x"bf",x"97",x"eb",x"ce"),
   364 => (x"e2",x"d6",x"c2",x"48"),
   365 => (x"48",x"4c",x"70",x"58"),
   366 => (x"d6",x"c2",x"88",x"c1"),
   367 => (x"ce",x"c2",x"58",x"e6"),
   368 => (x"49",x"bf",x"97",x"ec"),
   369 => (x"ce",x"c2",x"81",x"75"),
   370 => (x"4a",x"bf",x"97",x"ed"),
   371 => (x"a1",x"72",x"32",x"c8"),
   372 => (x"f3",x"da",x"c2",x"7e"),
   373 => (x"c2",x"78",x"6e",x"48"),
   374 => (x"bf",x"97",x"ee",x"ce"),
   375 => (x"58",x"a6",x"c8",x"48"),
   376 => (x"bf",x"e6",x"d6",x"c2"),
   377 => (x"87",x"d4",x"c2",x"02"),
   378 => (x"bf",x"e5",x"ed",x"c0"),
   379 => (x"f0",x"cf",x"c2",x"49"),
   380 => (x"4b",x"c8",x"71",x"4a"),
   381 => (x"70",x"87",x"f3",x"e9"),
   382 => (x"c5",x"c0",x"02",x"98"),
   383 => (x"c3",x"48",x"c0",x"87"),
   384 => (x"d6",x"c2",x"87",x"f8"),
   385 => (x"c2",x"4c",x"bf",x"de"),
   386 => (x"c2",x"5c",x"c7",x"db"),
   387 => (x"bf",x"97",x"c3",x"cf"),
   388 => (x"c2",x"31",x"c8",x"49"),
   389 => (x"bf",x"97",x"c2",x"cf"),
   390 => (x"c2",x"49",x"a1",x"4a"),
   391 => (x"bf",x"97",x"c4",x"cf"),
   392 => (x"72",x"32",x"d0",x"4a"),
   393 => (x"cf",x"c2",x"49",x"a1"),
   394 => (x"4a",x"bf",x"97",x"c5"),
   395 => (x"a1",x"72",x"32",x"d8"),
   396 => (x"91",x"66",x"c4",x"49"),
   397 => (x"bf",x"f3",x"da",x"c2"),
   398 => (x"fb",x"da",x"c2",x"81"),
   399 => (x"cb",x"cf",x"c2",x"59"),
   400 => (x"c8",x"4a",x"bf",x"97"),
   401 => (x"ca",x"cf",x"c2",x"32"),
   402 => (x"a2",x"4b",x"bf",x"97"),
   403 => (x"cc",x"cf",x"c2",x"4a"),
   404 => (x"d0",x"4b",x"bf",x"97"),
   405 => (x"4a",x"a2",x"73",x"33"),
   406 => (x"97",x"cd",x"cf",x"c2"),
   407 => (x"9b",x"cf",x"4b",x"bf"),
   408 => (x"a2",x"73",x"33",x"d8"),
   409 => (x"ff",x"da",x"c2",x"4a"),
   410 => (x"fb",x"da",x"c2",x"5a"),
   411 => (x"8a",x"c2",x"4a",x"bf"),
   412 => (x"da",x"c2",x"92",x"74"),
   413 => (x"a1",x"72",x"48",x"ff"),
   414 => (x"87",x"ca",x"c1",x"78"),
   415 => (x"97",x"f0",x"ce",x"c2"),
   416 => (x"31",x"c8",x"49",x"bf"),
   417 => (x"97",x"ef",x"ce",x"c2"),
   418 => (x"49",x"a1",x"4a",x"bf"),
   419 => (x"59",x"ee",x"d6",x"c2"),
   420 => (x"bf",x"ea",x"d6",x"c2"),
   421 => (x"c7",x"31",x"c5",x"49"),
   422 => (x"29",x"c9",x"81",x"ff"),
   423 => (x"59",x"c7",x"db",x"c2"),
   424 => (x"97",x"f5",x"ce",x"c2"),
   425 => (x"32",x"c8",x"4a",x"bf"),
   426 => (x"97",x"f4",x"ce",x"c2"),
   427 => (x"4a",x"a2",x"4b",x"bf"),
   428 => (x"6e",x"92",x"66",x"c4"),
   429 => (x"c3",x"db",x"c2",x"82"),
   430 => (x"fb",x"da",x"c2",x"5a"),
   431 => (x"c2",x"78",x"c0",x"48"),
   432 => (x"72",x"48",x"f7",x"da"),
   433 => (x"db",x"c2",x"78",x"a1"),
   434 => (x"da",x"c2",x"48",x"c7"),
   435 => (x"c2",x"78",x"bf",x"fb"),
   436 => (x"c2",x"48",x"cb",x"db"),
   437 => (x"78",x"bf",x"ff",x"da"),
   438 => (x"bf",x"e6",x"d6",x"c2"),
   439 => (x"87",x"c9",x"c0",x"02"),
   440 => (x"30",x"c4",x"48",x"74"),
   441 => (x"c9",x"c0",x"7e",x"70"),
   442 => (x"c3",x"db",x"c2",x"87"),
   443 => (x"30",x"c4",x"48",x"bf"),
   444 => (x"d6",x"c2",x"7e",x"70"),
   445 => (x"78",x"6e",x"48",x"ea"),
   446 => (x"8e",x"f8",x"48",x"c1"),
   447 => (x"4c",x"26",x"4d",x"26"),
   448 => (x"4f",x"26",x"4b",x"26"),
   449 => (x"5c",x"5b",x"5e",x"0e"),
   450 => (x"4a",x"71",x"0e",x"5d"),
   451 => (x"bf",x"e6",x"d6",x"c2"),
   452 => (x"72",x"87",x"cb",x"02"),
   453 => (x"72",x"2b",x"c7",x"4b"),
   454 => (x"9c",x"ff",x"c1",x"4c"),
   455 => (x"4b",x"72",x"87",x"c9"),
   456 => (x"4c",x"72",x"2b",x"c8"),
   457 => (x"c2",x"9c",x"ff",x"c3"),
   458 => (x"83",x"bf",x"f3",x"da"),
   459 => (x"bf",x"e1",x"ed",x"c0"),
   460 => (x"87",x"d9",x"02",x"ab"),
   461 => (x"5b",x"e5",x"ed",x"c0"),
   462 => (x"1e",x"de",x"ce",x"c2"),
   463 => (x"fd",x"f0",x"49",x"73"),
   464 => (x"70",x"86",x"c4",x"87"),
   465 => (x"87",x"c5",x"05",x"98"),
   466 => (x"e6",x"c0",x"48",x"c0"),
   467 => (x"e6",x"d6",x"c2",x"87"),
   468 => (x"87",x"d2",x"02",x"bf"),
   469 => (x"91",x"c4",x"49",x"74"),
   470 => (x"81",x"de",x"ce",x"c2"),
   471 => (x"ff",x"cf",x"4d",x"69"),
   472 => (x"9d",x"ff",x"ff",x"ff"),
   473 => (x"49",x"74",x"87",x"cb"),
   474 => (x"ce",x"c2",x"91",x"c2"),
   475 => (x"69",x"9f",x"81",x"de"),
   476 => (x"fe",x"48",x"75",x"4d"),
   477 => (x"5e",x"0e",x"87",x"c6"),
   478 => (x"0e",x"5d",x"5c",x"5b"),
   479 => (x"c0",x"4d",x"71",x"1e"),
   480 => (x"c8",x"49",x"c1",x"1e"),
   481 => (x"86",x"c4",x"87",x"c4"),
   482 => (x"02",x"9c",x"4c",x"70"),
   483 => (x"c2",x"87",x"c0",x"c1"),
   484 => (x"75",x"4a",x"ee",x"d6"),
   485 => (x"87",x"f7",x"e2",x"49"),
   486 => (x"c0",x"02",x"98",x"70"),
   487 => (x"4a",x"74",x"87",x"f1"),
   488 => (x"4b",x"cb",x"49",x"75"),
   489 => (x"70",x"87",x"dd",x"e3"),
   490 => (x"e2",x"c0",x"02",x"98"),
   491 => (x"74",x"1e",x"c0",x"87"),
   492 => (x"87",x"c7",x"02",x"9c"),
   493 => (x"c0",x"48",x"a6",x"c4"),
   494 => (x"c4",x"87",x"c5",x"78"),
   495 => (x"78",x"c1",x"48",x"a6"),
   496 => (x"c7",x"49",x"66",x"c4"),
   497 => (x"86",x"c4",x"87",x"c4"),
   498 => (x"05",x"9c",x"4c",x"70"),
   499 => (x"74",x"87",x"c0",x"ff"),
   500 => (x"e7",x"fc",x"26",x"48"),
   501 => (x"5b",x"5e",x"0e",x"87"),
   502 => (x"1e",x"0e",x"5d",x"5c"),
   503 => (x"05",x"9b",x"4b",x"71"),
   504 => (x"48",x"c0",x"87",x"c5"),
   505 => (x"c8",x"87",x"e5",x"c1"),
   506 => (x"7d",x"c0",x"4d",x"a3"),
   507 => (x"c7",x"02",x"66",x"d4"),
   508 => (x"97",x"66",x"d4",x"87"),
   509 => (x"87",x"c5",x"05",x"bf"),
   510 => (x"cf",x"c1",x"48",x"c0"),
   511 => (x"49",x"66",x"d4",x"87"),
   512 => (x"70",x"87",x"f3",x"fd"),
   513 => (x"c1",x"02",x"9c",x"4c"),
   514 => (x"a4",x"dc",x"87",x"c0"),
   515 => (x"da",x"7d",x"69",x"49"),
   516 => (x"a3",x"c4",x"49",x"a4"),
   517 => (x"7a",x"69",x"9f",x"4a"),
   518 => (x"bf",x"e6",x"d6",x"c2"),
   519 => (x"d4",x"87",x"d2",x"02"),
   520 => (x"69",x"9f",x"49",x"a4"),
   521 => (x"ff",x"ff",x"c0",x"49"),
   522 => (x"d0",x"48",x"71",x"99"),
   523 => (x"c2",x"7e",x"70",x"30"),
   524 => (x"6e",x"7e",x"c0",x"87"),
   525 => (x"80",x"6a",x"48",x"49"),
   526 => (x"7b",x"c0",x"7a",x"70"),
   527 => (x"6a",x"49",x"a3",x"cc"),
   528 => (x"49",x"a3",x"d0",x"79"),
   529 => (x"48",x"74",x"79",x"c0"),
   530 => (x"48",x"c0",x"87",x"c2"),
   531 => (x"87",x"ec",x"fa",x"26"),
   532 => (x"5c",x"5b",x"5e",x"0e"),
   533 => (x"4c",x"71",x"0e",x"5d"),
   534 => (x"48",x"e1",x"ed",x"c0"),
   535 => (x"9c",x"74",x"78",x"ff"),
   536 => (x"87",x"ca",x"c1",x"02"),
   537 => (x"69",x"49",x"a4",x"c8"),
   538 => (x"87",x"c2",x"c1",x"02"),
   539 => (x"6c",x"4a",x"66",x"d0"),
   540 => (x"a6",x"d4",x"82",x"49"),
   541 => (x"4d",x"66",x"d0",x"5a"),
   542 => (x"e2",x"d6",x"c2",x"b9"),
   543 => (x"ba",x"ff",x"4a",x"bf"),
   544 => (x"99",x"71",x"99",x"72"),
   545 => (x"87",x"e4",x"c0",x"02"),
   546 => (x"6b",x"4b",x"a4",x"c4"),
   547 => (x"87",x"f4",x"f9",x"49"),
   548 => (x"d6",x"c2",x"7b",x"70"),
   549 => (x"6c",x"49",x"bf",x"de"),
   550 => (x"75",x"7c",x"71",x"81"),
   551 => (x"e2",x"d6",x"c2",x"b9"),
   552 => (x"ba",x"ff",x"4a",x"bf"),
   553 => (x"99",x"71",x"99",x"72"),
   554 => (x"87",x"dc",x"ff",x"05"),
   555 => (x"cb",x"f9",x"7c",x"75"),
   556 => (x"1e",x"73",x"1e",x"87"),
   557 => (x"02",x"9b",x"4b",x"71"),
   558 => (x"a3",x"c8",x"87",x"c7"),
   559 => (x"c5",x"05",x"69",x"49"),
   560 => (x"c0",x"48",x"c0",x"87"),
   561 => (x"da",x"c2",x"87",x"eb"),
   562 => (x"c4",x"4a",x"bf",x"f7"),
   563 => (x"49",x"69",x"49",x"a3"),
   564 => (x"d6",x"c2",x"89",x"c2"),
   565 => (x"71",x"91",x"bf",x"de"),
   566 => (x"d6",x"c2",x"4a",x"a2"),
   567 => (x"6b",x"49",x"bf",x"e2"),
   568 => (x"4a",x"a2",x"71",x"99"),
   569 => (x"72",x"1e",x"66",x"c8"),
   570 => (x"87",x"d2",x"ea",x"49"),
   571 => (x"49",x"70",x"86",x"c4"),
   572 => (x"87",x"cc",x"f8",x"48"),
   573 => (x"71",x"1e",x"73",x"1e"),
   574 => (x"c0",x"02",x"9b",x"4b"),
   575 => (x"db",x"c2",x"87",x"e4"),
   576 => (x"4a",x"73",x"5b",x"cb"),
   577 => (x"d6",x"c2",x"8a",x"c2"),
   578 => (x"92",x"49",x"bf",x"de"),
   579 => (x"bf",x"f7",x"da",x"c2"),
   580 => (x"c2",x"80",x"72",x"48"),
   581 => (x"71",x"58",x"cf",x"db"),
   582 => (x"c2",x"30",x"c4",x"48"),
   583 => (x"c0",x"58",x"ee",x"d6"),
   584 => (x"db",x"c2",x"87",x"ed"),
   585 => (x"da",x"c2",x"48",x"c7"),
   586 => (x"c2",x"78",x"bf",x"fb"),
   587 => (x"c2",x"48",x"cb",x"db"),
   588 => (x"78",x"bf",x"ff",x"da"),
   589 => (x"bf",x"e6",x"d6",x"c2"),
   590 => (x"c2",x"87",x"c9",x"02"),
   591 => (x"49",x"bf",x"de",x"d6"),
   592 => (x"87",x"c7",x"31",x"c4"),
   593 => (x"bf",x"c3",x"db",x"c2"),
   594 => (x"c2",x"31",x"c4",x"49"),
   595 => (x"f6",x"59",x"ee",x"d6"),
   596 => (x"5e",x"0e",x"87",x"ee"),
   597 => (x"71",x"0e",x"5c",x"5b"),
   598 => (x"72",x"4b",x"c0",x"4a"),
   599 => (x"e1",x"c0",x"02",x"9a"),
   600 => (x"49",x"a2",x"da",x"87"),
   601 => (x"c2",x"4b",x"69",x"9f"),
   602 => (x"02",x"bf",x"e6",x"d6"),
   603 => (x"a2",x"d4",x"87",x"cf"),
   604 => (x"49",x"69",x"9f",x"49"),
   605 => (x"ff",x"ff",x"c0",x"4c"),
   606 => (x"c2",x"34",x"d0",x"9c"),
   607 => (x"74",x"4c",x"c0",x"87"),
   608 => (x"49",x"73",x"b3",x"49"),
   609 => (x"f5",x"87",x"ed",x"fd"),
   610 => (x"5e",x"0e",x"87",x"f4"),
   611 => (x"0e",x"5d",x"5c",x"5b"),
   612 => (x"4a",x"71",x"86",x"f4"),
   613 => (x"9a",x"72",x"7e",x"c0"),
   614 => (x"c2",x"87",x"d8",x"02"),
   615 => (x"c0",x"48",x"da",x"ce"),
   616 => (x"d2",x"ce",x"c2",x"78"),
   617 => (x"cb",x"db",x"c2",x"48"),
   618 => (x"ce",x"c2",x"78",x"bf"),
   619 => (x"db",x"c2",x"48",x"d6"),
   620 => (x"c2",x"78",x"bf",x"c7"),
   621 => (x"c0",x"48",x"fb",x"d6"),
   622 => (x"ea",x"d6",x"c2",x"50"),
   623 => (x"ce",x"c2",x"49",x"bf"),
   624 => (x"71",x"4a",x"bf",x"da"),
   625 => (x"ff",x"c3",x"03",x"aa"),
   626 => (x"cf",x"49",x"72",x"87"),
   627 => (x"e0",x"c0",x"05",x"99"),
   628 => (x"de",x"ce",x"c2",x"87"),
   629 => (x"d2",x"ce",x"c2",x"1e"),
   630 => (x"ce",x"c2",x"49",x"bf"),
   631 => (x"a1",x"c1",x"48",x"d2"),
   632 => (x"d9",x"e6",x"71",x"78"),
   633 => (x"c0",x"86",x"c4",x"87"),
   634 => (x"c2",x"48",x"dd",x"ed"),
   635 => (x"cc",x"78",x"de",x"ce"),
   636 => (x"dd",x"ed",x"c0",x"87"),
   637 => (x"e0",x"c0",x"48",x"bf"),
   638 => (x"e1",x"ed",x"c0",x"80"),
   639 => (x"da",x"ce",x"c2",x"58"),
   640 => (x"80",x"c1",x"48",x"bf"),
   641 => (x"58",x"de",x"ce",x"c2"),
   642 => (x"00",x"0b",x"5d",x"27"),
   643 => (x"bf",x"97",x"bf",x"00"),
   644 => (x"c2",x"02",x"9d",x"4d"),
   645 => (x"e5",x"c3",x"87",x"e2"),
   646 => (x"db",x"c2",x"02",x"ad"),
   647 => (x"dd",x"ed",x"c0",x"87"),
   648 => (x"a3",x"cb",x"4b",x"bf"),
   649 => (x"cf",x"4c",x"11",x"49"),
   650 => (x"d2",x"c1",x"05",x"ac"),
   651 => (x"df",x"49",x"75",x"87"),
   652 => (x"cd",x"89",x"c1",x"99"),
   653 => (x"ee",x"d6",x"c2",x"91"),
   654 => (x"4a",x"a3",x"c1",x"81"),
   655 => (x"a3",x"c3",x"51",x"12"),
   656 => (x"c5",x"51",x"12",x"4a"),
   657 => (x"51",x"12",x"4a",x"a3"),
   658 => (x"12",x"4a",x"a3",x"c7"),
   659 => (x"4a",x"a3",x"c9",x"51"),
   660 => (x"a3",x"ce",x"51",x"12"),
   661 => (x"d0",x"51",x"12",x"4a"),
   662 => (x"51",x"12",x"4a",x"a3"),
   663 => (x"12",x"4a",x"a3",x"d2"),
   664 => (x"4a",x"a3",x"d4",x"51"),
   665 => (x"a3",x"d6",x"51",x"12"),
   666 => (x"d8",x"51",x"12",x"4a"),
   667 => (x"51",x"12",x"4a",x"a3"),
   668 => (x"12",x"4a",x"a3",x"dc"),
   669 => (x"4a",x"a3",x"de",x"51"),
   670 => (x"7e",x"c1",x"51",x"12"),
   671 => (x"74",x"87",x"f9",x"c0"),
   672 => (x"05",x"99",x"c8",x"49"),
   673 => (x"74",x"87",x"ea",x"c0"),
   674 => (x"05",x"99",x"d0",x"49"),
   675 => (x"66",x"dc",x"87",x"d0"),
   676 => (x"87",x"ca",x"c0",x"02"),
   677 => (x"66",x"dc",x"49",x"73"),
   678 => (x"02",x"98",x"70",x"0f"),
   679 => (x"05",x"6e",x"87",x"d3"),
   680 => (x"c2",x"87",x"c6",x"c0"),
   681 => (x"c0",x"48",x"ee",x"d6"),
   682 => (x"dd",x"ed",x"c0",x"50"),
   683 => (x"e7",x"c2",x"48",x"bf"),
   684 => (x"fb",x"d6",x"c2",x"87"),
   685 => (x"7e",x"50",x"c0",x"48"),
   686 => (x"bf",x"ea",x"d6",x"c2"),
   687 => (x"da",x"ce",x"c2",x"49"),
   688 => (x"aa",x"71",x"4a",x"bf"),
   689 => (x"87",x"c1",x"fc",x"04"),
   690 => (x"bf",x"cb",x"db",x"c2"),
   691 => (x"87",x"c8",x"c0",x"05"),
   692 => (x"bf",x"e6",x"d6",x"c2"),
   693 => (x"87",x"fe",x"c1",x"02"),
   694 => (x"48",x"e1",x"ed",x"c0"),
   695 => (x"ce",x"c2",x"78",x"ff"),
   696 => (x"f0",x"49",x"bf",x"d6"),
   697 => (x"49",x"70",x"87",x"de"),
   698 => (x"59",x"da",x"ce",x"c2"),
   699 => (x"c2",x"48",x"a6",x"c4"),
   700 => (x"78",x"bf",x"d6",x"ce"),
   701 => (x"bf",x"e6",x"d6",x"c2"),
   702 => (x"87",x"d8",x"c0",x"02"),
   703 => (x"cf",x"49",x"66",x"c4"),
   704 => (x"f8",x"ff",x"ff",x"ff"),
   705 => (x"c0",x"02",x"a9",x"99"),
   706 => (x"4d",x"c0",x"87",x"c5"),
   707 => (x"c1",x"87",x"e1",x"c0"),
   708 => (x"87",x"dc",x"c0",x"4d"),
   709 => (x"cf",x"49",x"66",x"c4"),
   710 => (x"a9",x"99",x"f8",x"ff"),
   711 => (x"87",x"c8",x"c0",x"02"),
   712 => (x"c0",x"48",x"a6",x"c8"),
   713 => (x"87",x"c5",x"c0",x"78"),
   714 => (x"c1",x"48",x"a6",x"c8"),
   715 => (x"4d",x"66",x"c8",x"78"),
   716 => (x"c0",x"05",x"9d",x"75"),
   717 => (x"66",x"c4",x"87",x"e0"),
   718 => (x"c2",x"89",x"c2",x"49"),
   719 => (x"4a",x"bf",x"de",x"d6"),
   720 => (x"f7",x"da",x"c2",x"91"),
   721 => (x"ce",x"c2",x"4a",x"bf"),
   722 => (x"a1",x"72",x"48",x"d2"),
   723 => (x"da",x"ce",x"c2",x"78"),
   724 => (x"f9",x"78",x"c0",x"48"),
   725 => (x"48",x"c0",x"87",x"e3"),
   726 => (x"df",x"ee",x"8e",x"f4"),
   727 => (x"00",x"00",x"00",x"87"),
   728 => (x"ff",x"ff",x"ff",x"00"),
   729 => (x"00",x"0b",x"6d",x"ff"),
   730 => (x"00",x"0b",x"76",x"00"),
   731 => (x"54",x"41",x"46",x"00"),
   732 => (x"20",x"20",x"32",x"33"),
   733 => (x"41",x"46",x"00",x"20"),
   734 => (x"20",x"36",x"31",x"54"),
   735 => (x"1e",x"00",x"20",x"20"),
   736 => (x"c3",x"48",x"d4",x"ff"),
   737 => (x"48",x"68",x"78",x"ff"),
   738 => (x"ff",x"1e",x"4f",x"26"),
   739 => (x"ff",x"c3",x"48",x"d4"),
   740 => (x"48",x"d0",x"ff",x"78"),
   741 => (x"ff",x"78",x"e1",x"c8"),
   742 => (x"78",x"d4",x"48",x"d4"),
   743 => (x"48",x"cf",x"db",x"c2"),
   744 => (x"50",x"bf",x"d4",x"ff"),
   745 => (x"ff",x"1e",x"4f",x"26"),
   746 => (x"e0",x"c0",x"48",x"d0"),
   747 => (x"1e",x"4f",x"26",x"78"),
   748 => (x"70",x"87",x"cc",x"ff"),
   749 => (x"c6",x"02",x"99",x"49"),
   750 => (x"a9",x"fb",x"c0",x"87"),
   751 => (x"71",x"87",x"f1",x"05"),
   752 => (x"0e",x"4f",x"26",x"48"),
   753 => (x"0e",x"5c",x"5b",x"5e"),
   754 => (x"4c",x"c0",x"4b",x"71"),
   755 => (x"70",x"87",x"f0",x"fe"),
   756 => (x"c0",x"02",x"99",x"49"),
   757 => (x"ec",x"c0",x"87",x"f9"),
   758 => (x"f2",x"c0",x"02",x"a9"),
   759 => (x"a9",x"fb",x"c0",x"87"),
   760 => (x"87",x"eb",x"c0",x"02"),
   761 => (x"ac",x"b7",x"66",x"cc"),
   762 => (x"d0",x"87",x"c7",x"03"),
   763 => (x"87",x"c2",x"02",x"66"),
   764 => (x"99",x"71",x"53",x"71"),
   765 => (x"c1",x"87",x"c2",x"02"),
   766 => (x"87",x"c3",x"fe",x"84"),
   767 => (x"02",x"99",x"49",x"70"),
   768 => (x"ec",x"c0",x"87",x"cd"),
   769 => (x"87",x"c7",x"02",x"a9"),
   770 => (x"05",x"a9",x"fb",x"c0"),
   771 => (x"d0",x"87",x"d5",x"ff"),
   772 => (x"87",x"c3",x"02",x"66"),
   773 => (x"c0",x"7b",x"97",x"c0"),
   774 => (x"c4",x"05",x"a9",x"ec"),
   775 => (x"c5",x"4a",x"74",x"87"),
   776 => (x"c0",x"4a",x"74",x"87"),
   777 => (x"48",x"72",x"8a",x"0a"),
   778 => (x"4d",x"26",x"87",x"c2"),
   779 => (x"4b",x"26",x"4c",x"26"),
   780 => (x"fd",x"1e",x"4f",x"26"),
   781 => (x"49",x"70",x"87",x"c9"),
   782 => (x"a9",x"b7",x"f0",x"c0"),
   783 => (x"c0",x"87",x"ca",x"04"),
   784 => (x"01",x"a9",x"b7",x"f9"),
   785 => (x"f0",x"c0",x"87",x"c3"),
   786 => (x"b7",x"c1",x"c1",x"89"),
   787 => (x"87",x"ca",x"04",x"a9"),
   788 => (x"a9",x"b7",x"da",x"c1"),
   789 => (x"c0",x"87",x"c3",x"01"),
   790 => (x"48",x"71",x"89",x"f7"),
   791 => (x"5e",x"0e",x"4f",x"26"),
   792 => (x"71",x"0e",x"5c",x"5b"),
   793 => (x"4c",x"d4",x"ff",x"4a"),
   794 => (x"ea",x"c0",x"49",x"72"),
   795 => (x"9b",x"4b",x"70",x"87"),
   796 => (x"c1",x"87",x"c2",x"02"),
   797 => (x"48",x"d0",x"ff",x"8b"),
   798 => (x"c1",x"78",x"c5",x"c8"),
   799 => (x"49",x"73",x"7c",x"d5"),
   800 => (x"cd",x"c2",x"31",x"c6"),
   801 => (x"4a",x"bf",x"97",x"ca"),
   802 => (x"70",x"b0",x"71",x"48"),
   803 => (x"48",x"d0",x"ff",x"7c"),
   804 => (x"48",x"73",x"78",x"c4"),
   805 => (x"0e",x"87",x"d5",x"fe"),
   806 => (x"5d",x"5c",x"5b",x"5e"),
   807 => (x"71",x"86",x"f8",x"0e"),
   808 => (x"fb",x"7e",x"c0",x"4c"),
   809 => (x"4b",x"c0",x"87",x"e4"),
   810 => (x"97",x"c4",x"f5",x"c0"),
   811 => (x"a9",x"c0",x"49",x"bf"),
   812 => (x"fb",x"87",x"cf",x"04"),
   813 => (x"83",x"c1",x"87",x"f9"),
   814 => (x"97",x"c4",x"f5",x"c0"),
   815 => (x"06",x"ab",x"49",x"bf"),
   816 => (x"f5",x"c0",x"87",x"f1"),
   817 => (x"02",x"bf",x"97",x"c4"),
   818 => (x"f2",x"fa",x"87",x"cf"),
   819 => (x"99",x"49",x"70",x"87"),
   820 => (x"c0",x"87",x"c6",x"02"),
   821 => (x"f1",x"05",x"a9",x"ec"),
   822 => (x"fa",x"4b",x"c0",x"87"),
   823 => (x"4d",x"70",x"87",x"e1"),
   824 => (x"c8",x"87",x"dc",x"fa"),
   825 => (x"d6",x"fa",x"58",x"a6"),
   826 => (x"c1",x"4a",x"70",x"87"),
   827 => (x"49",x"a4",x"c8",x"83"),
   828 => (x"ad",x"49",x"69",x"97"),
   829 => (x"c0",x"87",x"c7",x"02"),
   830 => (x"c0",x"05",x"ad",x"ff"),
   831 => (x"a4",x"c9",x"87",x"e7"),
   832 => (x"49",x"69",x"97",x"49"),
   833 => (x"02",x"a9",x"66",x"c4"),
   834 => (x"c0",x"48",x"87",x"c7"),
   835 => (x"d4",x"05",x"a8",x"ff"),
   836 => (x"49",x"a4",x"ca",x"87"),
   837 => (x"aa",x"49",x"69",x"97"),
   838 => (x"c0",x"87",x"c6",x"02"),
   839 => (x"c4",x"05",x"aa",x"ff"),
   840 => (x"d0",x"7e",x"c1",x"87"),
   841 => (x"ad",x"ec",x"c0",x"87"),
   842 => (x"c0",x"87",x"c6",x"02"),
   843 => (x"c4",x"05",x"ad",x"fb"),
   844 => (x"c1",x"4b",x"c0",x"87"),
   845 => (x"fe",x"02",x"6e",x"7e"),
   846 => (x"e9",x"f9",x"87",x"e1"),
   847 => (x"f8",x"48",x"73",x"87"),
   848 => (x"87",x"e6",x"fb",x"8e"),
   849 => (x"5b",x"5e",x"0e",x"00"),
   850 => (x"1e",x"0e",x"5d",x"5c"),
   851 => (x"4c",x"c0",x"4b",x"71"),
   852 => (x"c0",x"04",x"ab",x"4d"),
   853 => (x"f2",x"c0",x"87",x"e8"),
   854 => (x"9d",x"75",x"1e",x"d7"),
   855 => (x"c0",x"87",x"c4",x"02"),
   856 => (x"c1",x"87",x"c2",x"4a"),
   857 => (x"f0",x"49",x"72",x"4a"),
   858 => (x"86",x"c4",x"87",x"e0"),
   859 => (x"84",x"c1",x"7e",x"70"),
   860 => (x"87",x"c2",x"05",x"6e"),
   861 => (x"85",x"c1",x"4c",x"73"),
   862 => (x"ff",x"06",x"ac",x"73"),
   863 => (x"48",x"6e",x"87",x"d8"),
   864 => (x"26",x"4d",x"26",x"26"),
   865 => (x"26",x"4b",x"26",x"4c"),
   866 => (x"5b",x"5e",x"0e",x"4f"),
   867 => (x"1e",x"0e",x"5d",x"5c"),
   868 => (x"de",x"49",x"4c",x"71"),
   869 => (x"e9",x"db",x"c2",x"91"),
   870 => (x"97",x"85",x"71",x"4d"),
   871 => (x"dd",x"c1",x"02",x"6d"),
   872 => (x"d4",x"db",x"c2",x"87"),
   873 => (x"82",x"74",x"4a",x"bf"),
   874 => (x"d8",x"fe",x"49",x"72"),
   875 => (x"6e",x"7e",x"70",x"87"),
   876 => (x"87",x"f3",x"c0",x"02"),
   877 => (x"4b",x"dc",x"db",x"c2"),
   878 => (x"49",x"cb",x"4a",x"6e"),
   879 => (x"87",x"e8",x"cb",x"ff"),
   880 => (x"93",x"cb",x"4b",x"74"),
   881 => (x"83",x"ee",x"d8",x"c1"),
   882 => (x"f8",x"c0",x"83",x"c4"),
   883 => (x"49",x"74",x"7b",x"c2"),
   884 => (x"87",x"d8",x"c2",x"c1"),
   885 => (x"db",x"c2",x"7b",x"75"),
   886 => (x"49",x"bf",x"97",x"e8"),
   887 => (x"dc",x"db",x"c2",x"1e"),
   888 => (x"d6",x"d5",x"c1",x"49"),
   889 => (x"74",x"86",x"c4",x"87"),
   890 => (x"ff",x"c1",x"c1",x"49"),
   891 => (x"c1",x"49",x"c0",x"87"),
   892 => (x"c2",x"87",x"de",x"c3"),
   893 => (x"c0",x"48",x"d0",x"db"),
   894 => (x"dd",x"49",x"c1",x"78"),
   895 => (x"fd",x"26",x"87",x"cb"),
   896 => (x"6f",x"4c",x"87",x"ff"),
   897 => (x"6e",x"69",x"64",x"61"),
   898 => (x"2e",x"2e",x"2e",x"67"),
   899 => (x"5b",x"5e",x"0e",x"00"),
   900 => (x"4b",x"71",x"0e",x"5c"),
   901 => (x"d4",x"db",x"c2",x"4a"),
   902 => (x"49",x"72",x"82",x"bf"),
   903 => (x"70",x"87",x"e6",x"fc"),
   904 => (x"c4",x"02",x"9c",x"4c"),
   905 => (x"e9",x"ec",x"49",x"87"),
   906 => (x"d4",x"db",x"c2",x"87"),
   907 => (x"c1",x"78",x"c0",x"48"),
   908 => (x"87",x"d5",x"dc",x"49"),
   909 => (x"0e",x"87",x"cc",x"fd"),
   910 => (x"5d",x"5c",x"5b",x"5e"),
   911 => (x"c2",x"86",x"f4",x"0e"),
   912 => (x"c0",x"4d",x"de",x"ce"),
   913 => (x"48",x"a6",x"c4",x"4c"),
   914 => (x"db",x"c2",x"78",x"c0"),
   915 => (x"c0",x"49",x"bf",x"d4"),
   916 => (x"c1",x"c1",x"06",x"a9"),
   917 => (x"de",x"ce",x"c2",x"87"),
   918 => (x"c0",x"02",x"98",x"48"),
   919 => (x"f2",x"c0",x"87",x"f8"),
   920 => (x"66",x"c8",x"1e",x"d7"),
   921 => (x"c4",x"87",x"c7",x"02"),
   922 => (x"78",x"c0",x"48",x"a6"),
   923 => (x"a6",x"c4",x"87",x"c5"),
   924 => (x"c4",x"78",x"c1",x"48"),
   925 => (x"d1",x"ec",x"49",x"66"),
   926 => (x"70",x"86",x"c4",x"87"),
   927 => (x"c4",x"84",x"c1",x"4d"),
   928 => (x"80",x"c1",x"48",x"66"),
   929 => (x"c2",x"58",x"a6",x"c8"),
   930 => (x"49",x"bf",x"d4",x"db"),
   931 => (x"87",x"c6",x"03",x"ac"),
   932 => (x"ff",x"05",x"9d",x"75"),
   933 => (x"4c",x"c0",x"87",x"c8"),
   934 => (x"c3",x"02",x"9d",x"75"),
   935 => (x"f2",x"c0",x"87",x"e0"),
   936 => (x"66",x"c8",x"1e",x"d7"),
   937 => (x"cc",x"87",x"c7",x"02"),
   938 => (x"78",x"c0",x"48",x"a6"),
   939 => (x"a6",x"cc",x"87",x"c5"),
   940 => (x"cc",x"78",x"c1",x"48"),
   941 => (x"d1",x"eb",x"49",x"66"),
   942 => (x"70",x"86",x"c4",x"87"),
   943 => (x"c2",x"02",x"6e",x"7e"),
   944 => (x"49",x"6e",x"87",x"e9"),
   945 => (x"69",x"97",x"81",x"cb"),
   946 => (x"02",x"99",x"d0",x"49"),
   947 => (x"c0",x"87",x"d6",x"c1"),
   948 => (x"74",x"4a",x"cd",x"f8"),
   949 => (x"c1",x"91",x"cb",x"49"),
   950 => (x"72",x"81",x"ee",x"d8"),
   951 => (x"c3",x"81",x"c8",x"79"),
   952 => (x"49",x"74",x"51",x"ff"),
   953 => (x"db",x"c2",x"91",x"de"),
   954 => (x"85",x"71",x"4d",x"e9"),
   955 => (x"7d",x"97",x"c1",x"c2"),
   956 => (x"c0",x"49",x"a5",x"c1"),
   957 => (x"d6",x"c2",x"51",x"e0"),
   958 => (x"02",x"bf",x"97",x"ee"),
   959 => (x"84",x"c1",x"87",x"d2"),
   960 => (x"c2",x"4b",x"a5",x"c2"),
   961 => (x"db",x"4a",x"ee",x"d6"),
   962 => (x"db",x"c6",x"ff",x"49"),
   963 => (x"87",x"db",x"c1",x"87"),
   964 => (x"c0",x"49",x"a5",x"cd"),
   965 => (x"c2",x"84",x"c1",x"51"),
   966 => (x"4a",x"6e",x"4b",x"a5"),
   967 => (x"c6",x"ff",x"49",x"cb"),
   968 => (x"c6",x"c1",x"87",x"c6"),
   969 => (x"c9",x"f6",x"c0",x"87"),
   970 => (x"cb",x"49",x"74",x"4a"),
   971 => (x"ee",x"d8",x"c1",x"91"),
   972 => (x"c2",x"79",x"72",x"81"),
   973 => (x"bf",x"97",x"ee",x"d6"),
   974 => (x"74",x"87",x"d8",x"02"),
   975 => (x"c1",x"91",x"de",x"49"),
   976 => (x"e9",x"db",x"c2",x"84"),
   977 => (x"c2",x"83",x"71",x"4b"),
   978 => (x"dd",x"4a",x"ee",x"d6"),
   979 => (x"d7",x"c5",x"ff",x"49"),
   980 => (x"74",x"87",x"d8",x"87"),
   981 => (x"c2",x"93",x"de",x"4b"),
   982 => (x"cb",x"83",x"e9",x"db"),
   983 => (x"51",x"c0",x"49",x"a3"),
   984 => (x"6e",x"73",x"84",x"c1"),
   985 => (x"ff",x"49",x"cb",x"4a"),
   986 => (x"c4",x"87",x"fd",x"c4"),
   987 => (x"80",x"c1",x"48",x"66"),
   988 => (x"c7",x"58",x"a6",x"c8"),
   989 => (x"c5",x"c0",x"03",x"ac"),
   990 => (x"fc",x"05",x"6e",x"87"),
   991 => (x"48",x"74",x"87",x"e0"),
   992 => (x"fc",x"f7",x"8e",x"f4"),
   993 => (x"1e",x"73",x"1e",x"87"),
   994 => (x"cb",x"49",x"4b",x"71"),
   995 => (x"ee",x"d8",x"c1",x"91"),
   996 => (x"4a",x"a1",x"c8",x"81"),
   997 => (x"48",x"ca",x"cd",x"c2"),
   998 => (x"a1",x"c9",x"50",x"12"),
   999 => (x"c4",x"f5",x"c0",x"4a"),
  1000 => (x"ca",x"50",x"12",x"48"),
  1001 => (x"e8",x"db",x"c2",x"81"),
  1002 => (x"c2",x"50",x"11",x"48"),
  1003 => (x"bf",x"97",x"e8",x"db"),
  1004 => (x"49",x"c0",x"1e",x"49"),
  1005 => (x"87",x"c3",x"ce",x"c1"),
  1006 => (x"48",x"d0",x"db",x"c2"),
  1007 => (x"49",x"c1",x"78",x"de"),
  1008 => (x"26",x"87",x"c6",x"d6"),
  1009 => (x"1e",x"87",x"fe",x"f6"),
  1010 => (x"cb",x"49",x"4a",x"71"),
  1011 => (x"ee",x"d8",x"c1",x"91"),
  1012 => (x"11",x"81",x"c8",x"81"),
  1013 => (x"d4",x"db",x"c2",x"48"),
  1014 => (x"d4",x"db",x"c2",x"58"),
  1015 => (x"c1",x"78",x"c0",x"48"),
  1016 => (x"87",x"e5",x"d5",x"49"),
  1017 => (x"c0",x"1e",x"4f",x"26"),
  1018 => (x"e4",x"fb",x"c0",x"49"),
  1019 => (x"1e",x"4f",x"26",x"87"),
  1020 => (x"d2",x"02",x"99",x"71"),
  1021 => (x"c3",x"da",x"c1",x"87"),
  1022 => (x"f7",x"50",x"c0",x"48"),
  1023 => (x"c7",x"ff",x"c0",x"80"),
  1024 => (x"e7",x"d8",x"c1",x"40"),
  1025 => (x"c1",x"87",x"ce",x"78"),
  1026 => (x"c1",x"48",x"ff",x"d9"),
  1027 => (x"fc",x"78",x"e0",x"d8"),
  1028 => (x"e6",x"ff",x"c0",x"80"),
  1029 => (x"0e",x"4f",x"26",x"78"),
  1030 => (x"0e",x"5c",x"5b",x"5e"),
  1031 => (x"cb",x"4a",x"4c",x"71"),
  1032 => (x"ee",x"d8",x"c1",x"92"),
  1033 => (x"49",x"a2",x"c8",x"82"),
  1034 => (x"97",x"4b",x"a2",x"c9"),
  1035 => (x"97",x"1e",x"4b",x"6b"),
  1036 => (x"ca",x"1e",x"49",x"69"),
  1037 => (x"c0",x"49",x"12",x"82"),
  1038 => (x"c0",x"87",x"df",x"e6"),
  1039 => (x"87",x"c9",x"d4",x"49"),
  1040 => (x"f8",x"c0",x"49",x"74"),
  1041 => (x"8e",x"f8",x"87",x"e6"),
  1042 => (x"1e",x"87",x"f8",x"f4"),
  1043 => (x"4b",x"71",x"1e",x"73"),
  1044 => (x"87",x"c3",x"ff",x"49"),
  1045 => (x"fe",x"fe",x"49",x"73"),
  1046 => (x"87",x"e9",x"f4",x"87"),
  1047 => (x"71",x"1e",x"73",x"1e"),
  1048 => (x"4a",x"a3",x"c6",x"4b"),
  1049 => (x"c1",x"87",x"db",x"02"),
  1050 => (x"87",x"d6",x"02",x"8a"),
  1051 => (x"da",x"c1",x"02",x"8a"),
  1052 => (x"c0",x"02",x"8a",x"87"),
  1053 => (x"02",x"8a",x"87",x"fc"),
  1054 => (x"8a",x"87",x"e1",x"c0"),
  1055 => (x"c1",x"87",x"cb",x"02"),
  1056 => (x"49",x"c7",x"87",x"db"),
  1057 => (x"c1",x"87",x"c0",x"fd"),
  1058 => (x"db",x"c2",x"87",x"de"),
  1059 => (x"c1",x"02",x"bf",x"d4"),
  1060 => (x"c1",x"48",x"87",x"cb"),
  1061 => (x"d8",x"db",x"c2",x"88"),
  1062 => (x"87",x"c1",x"c1",x"58"),
  1063 => (x"bf",x"d8",x"db",x"c2"),
  1064 => (x"87",x"f9",x"c0",x"02"),
  1065 => (x"bf",x"d4",x"db",x"c2"),
  1066 => (x"c2",x"80",x"c1",x"48"),
  1067 => (x"c0",x"58",x"d8",x"db"),
  1068 => (x"db",x"c2",x"87",x"eb"),
  1069 => (x"c6",x"49",x"bf",x"d4"),
  1070 => (x"d8",x"db",x"c2",x"89"),
  1071 => (x"a9",x"b7",x"c0",x"59"),
  1072 => (x"c2",x"87",x"da",x"03"),
  1073 => (x"c0",x"48",x"d4",x"db"),
  1074 => (x"c2",x"87",x"d2",x"78"),
  1075 => (x"02",x"bf",x"d8",x"db"),
  1076 => (x"db",x"c2",x"87",x"cb"),
  1077 => (x"c6",x"48",x"bf",x"d4"),
  1078 => (x"d8",x"db",x"c2",x"80"),
  1079 => (x"d1",x"49",x"c0",x"58"),
  1080 => (x"49",x"73",x"87",x"e7"),
  1081 => (x"87",x"c4",x"f6",x"c0"),
  1082 => (x"0e",x"87",x"da",x"f2"),
  1083 => (x"0e",x"5c",x"5b",x"5e"),
  1084 => (x"66",x"cc",x"4c",x"71"),
  1085 => (x"cb",x"4b",x"74",x"1e"),
  1086 => (x"ee",x"d8",x"c1",x"93"),
  1087 => (x"4a",x"a3",x"c4",x"83"),
  1088 => (x"fe",x"fe",x"49",x"6a"),
  1089 => (x"fe",x"c0",x"87",x"f2"),
  1090 => (x"a3",x"c8",x"7b",x"c5"),
  1091 => (x"51",x"66",x"d4",x"49"),
  1092 => (x"d8",x"49",x"a3",x"c9"),
  1093 => (x"a3",x"ca",x"51",x"66"),
  1094 => (x"51",x"66",x"dc",x"49"),
  1095 => (x"87",x"e3",x"f1",x"26"),
  1096 => (x"5c",x"5b",x"5e",x"0e"),
  1097 => (x"d0",x"ff",x"0e",x"5d"),
  1098 => (x"59",x"a6",x"d8",x"86"),
  1099 => (x"c0",x"48",x"a6",x"c4"),
  1100 => (x"c1",x"80",x"c4",x"78"),
  1101 => (x"c4",x"78",x"66",x"c4"),
  1102 => (x"c4",x"78",x"c1",x"80"),
  1103 => (x"c2",x"78",x"c1",x"80"),
  1104 => (x"c1",x"48",x"d8",x"db"),
  1105 => (x"d0",x"db",x"c2",x"78"),
  1106 => (x"a8",x"de",x"48",x"bf"),
  1107 => (x"f3",x"87",x"cb",x"05"),
  1108 => (x"49",x"70",x"87",x"e5"),
  1109 => (x"ce",x"59",x"a6",x"c8"),
  1110 => (x"ed",x"e8",x"87",x"f8"),
  1111 => (x"87",x"cf",x"e9",x"87"),
  1112 => (x"70",x"87",x"dc",x"e8"),
  1113 => (x"ac",x"fb",x"c0",x"4c"),
  1114 => (x"87",x"d0",x"c1",x"02"),
  1115 => (x"c1",x"05",x"66",x"d4"),
  1116 => (x"1e",x"c0",x"87",x"c2"),
  1117 => (x"c1",x"1e",x"c1",x"1e"),
  1118 => (x"c0",x"1e",x"e1",x"da"),
  1119 => (x"87",x"eb",x"fd",x"49"),
  1120 => (x"4a",x"66",x"d0",x"c1"),
  1121 => (x"49",x"6a",x"82",x"c4"),
  1122 => (x"51",x"74",x"81",x"c7"),
  1123 => (x"1e",x"d8",x"1e",x"c1"),
  1124 => (x"81",x"c8",x"49",x"6a"),
  1125 => (x"d8",x"87",x"ec",x"e8"),
  1126 => (x"66",x"c4",x"c1",x"86"),
  1127 => (x"01",x"a8",x"c0",x"48"),
  1128 => (x"a6",x"c4",x"87",x"c7"),
  1129 => (x"ce",x"78",x"c1",x"48"),
  1130 => (x"66",x"c4",x"c1",x"87"),
  1131 => (x"cc",x"88",x"c1",x"48"),
  1132 => (x"87",x"c3",x"58",x"a6"),
  1133 => (x"cc",x"87",x"f8",x"e7"),
  1134 => (x"78",x"c2",x"48",x"a6"),
  1135 => (x"cd",x"02",x"9c",x"74"),
  1136 => (x"66",x"c4",x"87",x"cc"),
  1137 => (x"66",x"c8",x"c1",x"48"),
  1138 => (x"c1",x"cd",x"03",x"a8"),
  1139 => (x"48",x"a6",x"d8",x"87"),
  1140 => (x"ea",x"e6",x"78",x"c0"),
  1141 => (x"c1",x"4c",x"70",x"87"),
  1142 => (x"c2",x"05",x"ac",x"d0"),
  1143 => (x"66",x"d8",x"87",x"d6"),
  1144 => (x"87",x"ce",x"e9",x"7e"),
  1145 => (x"a6",x"dc",x"49",x"70"),
  1146 => (x"87",x"d3",x"e6",x"59"),
  1147 => (x"ec",x"c0",x"4c",x"70"),
  1148 => (x"ea",x"c1",x"05",x"ac"),
  1149 => (x"49",x"66",x"c4",x"87"),
  1150 => (x"c0",x"c1",x"91",x"cb"),
  1151 => (x"a1",x"c4",x"81",x"66"),
  1152 => (x"c8",x"4d",x"6a",x"4a"),
  1153 => (x"66",x"d8",x"4a",x"a1"),
  1154 => (x"c7",x"ff",x"c0",x"52"),
  1155 => (x"87",x"ef",x"e5",x"79"),
  1156 => (x"02",x"9c",x"4c",x"70"),
  1157 => (x"fb",x"c0",x"87",x"d8"),
  1158 => (x"87",x"d2",x"02",x"ac"),
  1159 => (x"de",x"e5",x"55",x"74"),
  1160 => (x"9c",x"4c",x"70",x"87"),
  1161 => (x"c0",x"87",x"c7",x"02"),
  1162 => (x"ff",x"05",x"ac",x"fb"),
  1163 => (x"e0",x"c0",x"87",x"ee"),
  1164 => (x"55",x"c1",x"c2",x"55"),
  1165 => (x"d4",x"7d",x"97",x"c0"),
  1166 => (x"a9",x"6e",x"49",x"66"),
  1167 => (x"c4",x"87",x"db",x"05"),
  1168 => (x"66",x"c8",x"48",x"66"),
  1169 => (x"87",x"ca",x"04",x"a8"),
  1170 => (x"c1",x"48",x"66",x"c4"),
  1171 => (x"58",x"a6",x"c8",x"80"),
  1172 => (x"66",x"c8",x"87",x"c8"),
  1173 => (x"cc",x"88",x"c1",x"48"),
  1174 => (x"e2",x"e4",x"58",x"a6"),
  1175 => (x"c1",x"4c",x"70",x"87"),
  1176 => (x"c8",x"05",x"ac",x"d0"),
  1177 => (x"48",x"66",x"d0",x"87"),
  1178 => (x"a6",x"d4",x"80",x"c1"),
  1179 => (x"ac",x"d0",x"c1",x"58"),
  1180 => (x"87",x"ea",x"fd",x"02"),
  1181 => (x"d4",x"48",x"a6",x"dc"),
  1182 => (x"66",x"d8",x"78",x"66"),
  1183 => (x"a8",x"66",x"dc",x"48"),
  1184 => (x"87",x"dc",x"c9",x"05"),
  1185 => (x"48",x"a6",x"e0",x"c0"),
  1186 => (x"c4",x"78",x"f0",x"c0"),
  1187 => (x"78",x"66",x"cc",x"80"),
  1188 => (x"78",x"c0",x"80",x"c4"),
  1189 => (x"c0",x"48",x"74",x"7e"),
  1190 => (x"f0",x"c0",x"88",x"fb"),
  1191 => (x"98",x"70",x"58",x"a6"),
  1192 => (x"87",x"d7",x"c8",x"02"),
  1193 => (x"c0",x"88",x"cb",x"48"),
  1194 => (x"70",x"58",x"a6",x"f0"),
  1195 => (x"e9",x"c0",x"02",x"98"),
  1196 => (x"88",x"c9",x"48",x"87"),
  1197 => (x"58",x"a6",x"f0",x"c0"),
  1198 => (x"c3",x"02",x"98",x"70"),
  1199 => (x"c4",x"48",x"87",x"e1"),
  1200 => (x"a6",x"f0",x"c0",x"88"),
  1201 => (x"02",x"98",x"70",x"58"),
  1202 => (x"c1",x"48",x"87",x"d6"),
  1203 => (x"a6",x"f0",x"c0",x"88"),
  1204 => (x"02",x"98",x"70",x"58"),
  1205 => (x"c7",x"87",x"c8",x"c3"),
  1206 => (x"e0",x"c0",x"87",x"db"),
  1207 => (x"78",x"c0",x"48",x"a6"),
  1208 => (x"c1",x"48",x"66",x"cc"),
  1209 => (x"58",x"a6",x"d0",x"80"),
  1210 => (x"70",x"87",x"d4",x"e2"),
  1211 => (x"ac",x"ec",x"c0",x"4c"),
  1212 => (x"c0",x"87",x"d5",x"02"),
  1213 => (x"c6",x"02",x"66",x"e0"),
  1214 => (x"a6",x"e4",x"c0",x"87"),
  1215 => (x"74",x"87",x"c9",x"5c"),
  1216 => (x"88",x"f0",x"c0",x"48"),
  1217 => (x"58",x"a6",x"e8",x"c0"),
  1218 => (x"02",x"ac",x"ec",x"c0"),
  1219 => (x"ee",x"e1",x"87",x"cc"),
  1220 => (x"c0",x"4c",x"70",x"87"),
  1221 => (x"ff",x"05",x"ac",x"ec"),
  1222 => (x"e0",x"c0",x"87",x"f4"),
  1223 => (x"66",x"d4",x"1e",x"66"),
  1224 => (x"ec",x"c0",x"1e",x"49"),
  1225 => (x"da",x"c1",x"1e",x"66"),
  1226 => (x"66",x"d4",x"1e",x"e1"),
  1227 => (x"87",x"fb",x"f6",x"49"),
  1228 => (x"1e",x"ca",x"1e",x"c0"),
  1229 => (x"cb",x"49",x"66",x"dc"),
  1230 => (x"66",x"d8",x"c1",x"91"),
  1231 => (x"48",x"a6",x"d8",x"81"),
  1232 => (x"d8",x"78",x"a1",x"c4"),
  1233 => (x"e1",x"49",x"bf",x"66"),
  1234 => (x"86",x"d8",x"87",x"f9"),
  1235 => (x"06",x"a8",x"b7",x"c0"),
  1236 => (x"c1",x"87",x"c7",x"c1"),
  1237 => (x"c8",x"1e",x"de",x"1e"),
  1238 => (x"e1",x"49",x"bf",x"66"),
  1239 => (x"86",x"c8",x"87",x"e5"),
  1240 => (x"c0",x"48",x"49",x"70"),
  1241 => (x"e4",x"c0",x"88",x"08"),
  1242 => (x"b7",x"c0",x"58",x"a6"),
  1243 => (x"e9",x"c0",x"06",x"a8"),
  1244 => (x"66",x"e0",x"c0",x"87"),
  1245 => (x"a8",x"b7",x"dd",x"48"),
  1246 => (x"6e",x"87",x"df",x"03"),
  1247 => (x"e0",x"c0",x"49",x"bf"),
  1248 => (x"e0",x"c0",x"81",x"66"),
  1249 => (x"c1",x"49",x"66",x"51"),
  1250 => (x"81",x"bf",x"6e",x"81"),
  1251 => (x"c0",x"51",x"c1",x"c2"),
  1252 => (x"c2",x"49",x"66",x"e0"),
  1253 => (x"81",x"bf",x"6e",x"81"),
  1254 => (x"7e",x"c1",x"51",x"c0"),
  1255 => (x"e2",x"87",x"dc",x"c4"),
  1256 => (x"e4",x"c0",x"87",x"d0"),
  1257 => (x"c9",x"e2",x"58",x"a6"),
  1258 => (x"a6",x"e8",x"c0",x"87"),
  1259 => (x"a8",x"ec",x"c0",x"58"),
  1260 => (x"87",x"cb",x"c0",x"05"),
  1261 => (x"48",x"a6",x"e4",x"c0"),
  1262 => (x"78",x"66",x"e0",x"c0"),
  1263 => (x"ff",x"87",x"c4",x"c0"),
  1264 => (x"c4",x"87",x"fc",x"de"),
  1265 => (x"91",x"cb",x"49",x"66"),
  1266 => (x"48",x"66",x"c0",x"c1"),
  1267 => (x"7e",x"70",x"80",x"71"),
  1268 => (x"82",x"c8",x"4a",x"6e"),
  1269 => (x"81",x"ca",x"49",x"6e"),
  1270 => (x"51",x"66",x"e0",x"c0"),
  1271 => (x"49",x"66",x"e4",x"c0"),
  1272 => (x"e0",x"c0",x"81",x"c1"),
  1273 => (x"48",x"c1",x"89",x"66"),
  1274 => (x"49",x"70",x"30",x"71"),
  1275 => (x"97",x"71",x"89",x"c1"),
  1276 => (x"c5",x"df",x"c2",x"7a"),
  1277 => (x"e0",x"c0",x"49",x"bf"),
  1278 => (x"6a",x"97",x"29",x"66"),
  1279 => (x"98",x"71",x"48",x"4a"),
  1280 => (x"58",x"a6",x"f0",x"c0"),
  1281 => (x"81",x"c4",x"49",x"6e"),
  1282 => (x"66",x"dc",x"4d",x"69"),
  1283 => (x"a8",x"66",x"d8",x"48"),
  1284 => (x"87",x"c8",x"c0",x"02"),
  1285 => (x"c0",x"48",x"a6",x"d8"),
  1286 => (x"87",x"c5",x"c0",x"78"),
  1287 => (x"c1",x"48",x"a6",x"d8"),
  1288 => (x"1e",x"66",x"d8",x"78"),
  1289 => (x"75",x"1e",x"e0",x"c0"),
  1290 => (x"d6",x"de",x"ff",x"49"),
  1291 => (x"70",x"86",x"c8",x"87"),
  1292 => (x"ac",x"b7",x"c0",x"4c"),
  1293 => (x"87",x"d4",x"c1",x"06"),
  1294 => (x"e0",x"c0",x"85",x"74"),
  1295 => (x"75",x"89",x"74",x"49"),
  1296 => (x"c6",x"d5",x"c1",x"4b"),
  1297 => (x"f1",x"fe",x"71",x"4a"),
  1298 => (x"85",x"c2",x"87",x"de"),
  1299 => (x"48",x"66",x"e8",x"c0"),
  1300 => (x"ec",x"c0",x"80",x"c1"),
  1301 => (x"ec",x"c0",x"58",x"a6"),
  1302 => (x"81",x"c1",x"49",x"66"),
  1303 => (x"c0",x"02",x"a9",x"70"),
  1304 => (x"a6",x"d8",x"87",x"c8"),
  1305 => (x"c0",x"78",x"c0",x"48"),
  1306 => (x"a6",x"d8",x"87",x"c5"),
  1307 => (x"d8",x"78",x"c1",x"48"),
  1308 => (x"a4",x"c2",x"1e",x"66"),
  1309 => (x"48",x"e0",x"c0",x"49"),
  1310 => (x"49",x"70",x"88",x"71"),
  1311 => (x"ff",x"49",x"75",x"1e"),
  1312 => (x"c8",x"87",x"c0",x"dd"),
  1313 => (x"a8",x"b7",x"c0",x"86"),
  1314 => (x"87",x"c0",x"ff",x"01"),
  1315 => (x"02",x"66",x"e8",x"c0"),
  1316 => (x"6e",x"87",x"d1",x"c0"),
  1317 => (x"c0",x"81",x"c9",x"49"),
  1318 => (x"6e",x"51",x"66",x"e8"),
  1319 => (x"d7",x"c0",x"c1",x"48"),
  1320 => (x"87",x"cc",x"c0",x"78"),
  1321 => (x"81",x"c9",x"49",x"6e"),
  1322 => (x"48",x"6e",x"51",x"c2"),
  1323 => (x"78",x"cb",x"c1",x"c1"),
  1324 => (x"c6",x"c0",x"7e",x"c1"),
  1325 => (x"f6",x"db",x"ff",x"87"),
  1326 => (x"6e",x"4c",x"70",x"87"),
  1327 => (x"87",x"f5",x"c0",x"02"),
  1328 => (x"c8",x"48",x"66",x"c4"),
  1329 => (x"c0",x"04",x"a8",x"66"),
  1330 => (x"66",x"c4",x"87",x"cb"),
  1331 => (x"c8",x"80",x"c1",x"48"),
  1332 => (x"e0",x"c0",x"58",x"a6"),
  1333 => (x"48",x"66",x"c8",x"87"),
  1334 => (x"a6",x"cc",x"88",x"c1"),
  1335 => (x"87",x"d5",x"c0",x"58"),
  1336 => (x"05",x"ac",x"c6",x"c1"),
  1337 => (x"cc",x"87",x"c8",x"c0"),
  1338 => (x"80",x"c1",x"48",x"66"),
  1339 => (x"ff",x"58",x"a6",x"d0"),
  1340 => (x"70",x"87",x"fc",x"da"),
  1341 => (x"48",x"66",x"d0",x"4c"),
  1342 => (x"a6",x"d4",x"80",x"c1"),
  1343 => (x"02",x"9c",x"74",x"58"),
  1344 => (x"c4",x"87",x"cb",x"c0"),
  1345 => (x"c8",x"c1",x"48",x"66"),
  1346 => (x"f2",x"04",x"a8",x"66"),
  1347 => (x"da",x"ff",x"87",x"ff"),
  1348 => (x"66",x"c4",x"87",x"d4"),
  1349 => (x"03",x"a8",x"c7",x"48"),
  1350 => (x"c2",x"87",x"e5",x"c0"),
  1351 => (x"c0",x"48",x"d8",x"db"),
  1352 => (x"49",x"66",x"c4",x"78"),
  1353 => (x"c0",x"c1",x"91",x"cb"),
  1354 => (x"a1",x"c4",x"81",x"66"),
  1355 => (x"c0",x"4a",x"6a",x"4a"),
  1356 => (x"66",x"c4",x"79",x"52"),
  1357 => (x"c8",x"80",x"c1",x"48"),
  1358 => (x"a8",x"c7",x"58",x"a6"),
  1359 => (x"87",x"db",x"ff",x"04"),
  1360 => (x"e0",x"8e",x"d0",x"ff"),
  1361 => (x"20",x"3a",x"87",x"fb"),
  1362 => (x"1e",x"73",x"1e",x"00"),
  1363 => (x"02",x"9b",x"4b",x"71"),
  1364 => (x"db",x"c2",x"87",x"c6"),
  1365 => (x"78",x"c0",x"48",x"d4"),
  1366 => (x"db",x"c2",x"1e",x"c7"),
  1367 => (x"1e",x"49",x"bf",x"d4"),
  1368 => (x"1e",x"ee",x"d8",x"c1"),
  1369 => (x"bf",x"d0",x"db",x"c2"),
  1370 => (x"87",x"f4",x"ee",x"49"),
  1371 => (x"db",x"c2",x"86",x"cc"),
  1372 => (x"e9",x"49",x"bf",x"d0"),
  1373 => (x"9b",x"73",x"87",x"f9"),
  1374 => (x"c1",x"87",x"c8",x"02"),
  1375 => (x"c0",x"49",x"ee",x"d8"),
  1376 => (x"ff",x"87",x"fb",x"e4"),
  1377 => (x"1e",x"87",x"fe",x"df"),
  1378 => (x"48",x"ca",x"cd",x"c2"),
  1379 => (x"da",x"c1",x"50",x"c0"),
  1380 => (x"c0",x"49",x"bf",x"d1"),
  1381 => (x"c0",x"87",x"f7",x"f2"),
  1382 => (x"1e",x"4f",x"26",x"48"),
  1383 => (x"c1",x"87",x"e1",x"c7"),
  1384 => (x"87",x"e5",x"fe",x"49"),
  1385 => (x"87",x"fd",x"f3",x"fe"),
  1386 => (x"cd",x"02",x"98",x"70"),
  1387 => (x"d8",x"fb",x"fe",x"87"),
  1388 => (x"02",x"98",x"70",x"87"),
  1389 => (x"4a",x"c1",x"87",x"c4"),
  1390 => (x"4a",x"c0",x"87",x"c2"),
  1391 => (x"ce",x"05",x"9a",x"72"),
  1392 => (x"c1",x"1e",x"c0",x"87"),
  1393 => (x"c0",x"49",x"eb",x"d7"),
  1394 => (x"c4",x"87",x"c1",x"f0"),
  1395 => (x"c0",x"87",x"fe",x"86"),
  1396 => (x"f6",x"d7",x"c1",x"1e"),
  1397 => (x"f3",x"ef",x"c0",x"49"),
  1398 => (x"fe",x"1e",x"c0",x"87"),
  1399 => (x"49",x"70",x"87",x"e9"),
  1400 => (x"87",x"e8",x"ef",x"c0"),
  1401 => (x"f8",x"87",x"d8",x"c3"),
  1402 => (x"53",x"4f",x"26",x"8e"),
  1403 => (x"61",x"66",x"20",x"44"),
  1404 => (x"64",x"65",x"6c",x"69"),
  1405 => (x"6f",x"42",x"00",x"2e"),
  1406 => (x"6e",x"69",x"74",x"6f"),
  1407 => (x"2e",x"2e",x"2e",x"67"),
  1408 => (x"e7",x"c0",x"1e",x"00"),
  1409 => (x"87",x"fa",x"87",x"d4"),
  1410 => (x"c2",x"1e",x"4f",x"26"),
  1411 => (x"c0",x"48",x"d4",x"db"),
  1412 => (x"d0",x"db",x"c2",x"78"),
  1413 => (x"fe",x"78",x"c0",x"48"),
  1414 => (x"87",x"e5",x"87",x"c1"),
  1415 => (x"4f",x"26",x"48",x"c0"),
  1416 => (x"78",x"45",x"20",x"80"),
  1417 => (x"80",x"00",x"74",x"69"),
  1418 => (x"63",x"61",x"42",x"20"),
  1419 => (x"0f",x"c7",x"00",x"6b"),
  1420 => (x"26",x"e9",x"00",x"00"),
  1421 => (x"00",x"00",x"00",x"00"),
  1422 => (x"00",x"0f",x"c7",x"00"),
  1423 => (x"00",x"27",x"07",x"00"),
  1424 => (x"00",x"00",x"00",x"00"),
  1425 => (x"00",x"00",x"0f",x"c7"),
  1426 => (x"00",x"00",x"27",x"25"),
  1427 => (x"c7",x"00",x"00",x"00"),
  1428 => (x"43",x"00",x"00",x"0f"),
  1429 => (x"00",x"00",x"00",x"27"),
  1430 => (x"0f",x"c7",x"00",x"00"),
  1431 => (x"27",x"61",x"00",x"00"),
  1432 => (x"00",x"00",x"00",x"00"),
  1433 => (x"00",x"0f",x"c7",x"00"),
  1434 => (x"00",x"27",x"7f",x"00"),
  1435 => (x"00",x"00",x"00",x"00"),
  1436 => (x"00",x"00",x"0f",x"c7"),
  1437 => (x"00",x"00",x"27",x"9d"),
  1438 => (x"c7",x"00",x"00",x"00"),
  1439 => (x"00",x"00",x"00",x"0f"),
  1440 => (x"00",x"00",x"00",x"00"),
  1441 => (x"10",x"5c",x"00",x"00"),
  1442 => (x"00",x"00",x"00",x"00"),
  1443 => (x"00",x"00",x"00",x"00"),
  1444 => (x"00",x"16",x"95",x"00"),
  1445 => (x"4f",x"4f",x"42",x"00"),
  1446 => (x"20",x"20",x"20",x"54"),
  1447 => (x"4d",x"4f",x"52",x"20"),
  1448 => (x"61",x"6f",x"4c",x"00"),
  1449 => (x"2e",x"2a",x"20",x"64"),
  1450 => (x"f0",x"fe",x"1e",x"00"),
  1451 => (x"cd",x"78",x"c0",x"48"),
  1452 => (x"26",x"09",x"79",x"09"),
  1453 => (x"fe",x"1e",x"1e",x"4f"),
  1454 => (x"48",x"7e",x"bf",x"f0"),
  1455 => (x"1e",x"4f",x"26",x"26"),
  1456 => (x"c1",x"48",x"f0",x"fe"),
  1457 => (x"1e",x"4f",x"26",x"78"),
  1458 => (x"c0",x"48",x"f0",x"fe"),
  1459 => (x"1e",x"4f",x"26",x"78"),
  1460 => (x"52",x"c0",x"4a",x"71"),
  1461 => (x"0e",x"4f",x"26",x"52"),
  1462 => (x"5d",x"5c",x"5b",x"5e"),
  1463 => (x"71",x"86",x"f4",x"0e"),
  1464 => (x"7e",x"6d",x"97",x"4d"),
  1465 => (x"97",x"4c",x"a5",x"c1"),
  1466 => (x"a6",x"c8",x"48",x"6c"),
  1467 => (x"c4",x"48",x"6e",x"58"),
  1468 => (x"c5",x"05",x"a8",x"66"),
  1469 => (x"c0",x"48",x"ff",x"87"),
  1470 => (x"ca",x"ff",x"87",x"e6"),
  1471 => (x"49",x"a5",x"c2",x"87"),
  1472 => (x"71",x"4b",x"6c",x"97"),
  1473 => (x"6b",x"97",x"4b",x"a3"),
  1474 => (x"7e",x"6c",x"97",x"4b"),
  1475 => (x"80",x"c1",x"48",x"6e"),
  1476 => (x"c7",x"58",x"a6",x"c8"),
  1477 => (x"58",x"a6",x"cc",x"98"),
  1478 => (x"fe",x"7c",x"97",x"70"),
  1479 => (x"48",x"73",x"87",x"e1"),
  1480 => (x"4d",x"26",x"8e",x"f4"),
  1481 => (x"4b",x"26",x"4c",x"26"),
  1482 => (x"5e",x"0e",x"4f",x"26"),
  1483 => (x"f4",x"0e",x"5c",x"5b"),
  1484 => (x"d8",x"4c",x"71",x"86"),
  1485 => (x"ff",x"c3",x"4a",x"66"),
  1486 => (x"4b",x"a4",x"c2",x"9a"),
  1487 => (x"73",x"49",x"6c",x"97"),
  1488 => (x"51",x"72",x"49",x"a1"),
  1489 => (x"6e",x"7e",x"6c",x"97"),
  1490 => (x"c8",x"80",x"c1",x"48"),
  1491 => (x"98",x"c7",x"58",x"a6"),
  1492 => (x"70",x"58",x"a6",x"cc"),
  1493 => (x"ff",x"8e",x"f4",x"54"),
  1494 => (x"1e",x"1e",x"87",x"ca"),
  1495 => (x"e0",x"87",x"e8",x"fd"),
  1496 => (x"c0",x"49",x"4a",x"bf"),
  1497 => (x"02",x"99",x"c0",x"e0"),
  1498 => (x"1e",x"72",x"87",x"cb"),
  1499 => (x"49",x"fb",x"de",x"c2"),
  1500 => (x"c4",x"87",x"f7",x"fe"),
  1501 => (x"87",x"fd",x"fc",x"86"),
  1502 => (x"c2",x"fd",x"7e",x"70"),
  1503 => (x"4f",x"26",x"26",x"87"),
  1504 => (x"fb",x"de",x"c2",x"1e"),
  1505 => (x"87",x"c7",x"fd",x"49"),
  1506 => (x"49",x"da",x"dd",x"c1"),
  1507 => (x"c4",x"87",x"da",x"fc"),
  1508 => (x"4f",x"26",x"87",x"ff"),
  1509 => (x"5c",x"5b",x"5e",x"0e"),
  1510 => (x"df",x"c2",x"0e",x"5d"),
  1511 => (x"c1",x"4a",x"bf",x"da"),
  1512 => (x"49",x"bf",x"e8",x"df"),
  1513 => (x"71",x"bc",x"72",x"4c"),
  1514 => (x"87",x"db",x"fc",x"4d"),
  1515 => (x"49",x"74",x"4b",x"c0"),
  1516 => (x"d5",x"02",x"99",x"d0"),
  1517 => (x"d0",x"49",x"75",x"87"),
  1518 => (x"c0",x"1e",x"71",x"99"),
  1519 => (x"e0",x"e5",x"c1",x"1e"),
  1520 => (x"12",x"82",x"73",x"4a"),
  1521 => (x"87",x"e4",x"c0",x"49"),
  1522 => (x"2c",x"c1",x"86",x"c8"),
  1523 => (x"ab",x"c8",x"83",x"2d"),
  1524 => (x"87",x"da",x"ff",x"04"),
  1525 => (x"c1",x"87",x"e8",x"fb"),
  1526 => (x"c2",x"48",x"e8",x"df"),
  1527 => (x"78",x"bf",x"da",x"df"),
  1528 => (x"4c",x"26",x"4d",x"26"),
  1529 => (x"4f",x"26",x"4b",x"26"),
  1530 => (x"00",x"00",x"00",x"00"),
  1531 => (x"48",x"d0",x"ff",x"1e"),
  1532 => (x"ff",x"78",x"e1",x"c8"),
  1533 => (x"78",x"c5",x"48",x"d4"),
  1534 => (x"c3",x"02",x"66",x"c4"),
  1535 => (x"78",x"e0",x"c3",x"87"),
  1536 => (x"c6",x"02",x"66",x"c8"),
  1537 => (x"48",x"d4",x"ff",x"87"),
  1538 => (x"ff",x"78",x"f0",x"c3"),
  1539 => (x"78",x"71",x"48",x"d4"),
  1540 => (x"c8",x"48",x"d0",x"ff"),
  1541 => (x"e0",x"c0",x"78",x"e1"),
  1542 => (x"1e",x"4f",x"26",x"78"),
  1543 => (x"de",x"c2",x"1e",x"73"),
  1544 => (x"f2",x"fa",x"49",x"fb"),
  1545 => (x"c0",x"4a",x"70",x"87"),
  1546 => (x"c2",x"04",x"aa",x"b7"),
  1547 => (x"e0",x"c3",x"87",x"cd"),
  1548 => (x"87",x"c9",x"05",x"aa"),
  1549 => (x"48",x"c4",x"e3",x"c1"),
  1550 => (x"fe",x"c1",x"78",x"c1"),
  1551 => (x"aa",x"f0",x"c3",x"87"),
  1552 => (x"c1",x"87",x"c9",x"05"),
  1553 => (x"c1",x"48",x"c0",x"e3"),
  1554 => (x"87",x"df",x"c1",x"78"),
  1555 => (x"bf",x"c4",x"e3",x"c1"),
  1556 => (x"72",x"87",x"c7",x"02"),
  1557 => (x"b3",x"c0",x"c2",x"4b"),
  1558 => (x"4b",x"72",x"87",x"c2"),
  1559 => (x"bf",x"c0",x"e3",x"c1"),
  1560 => (x"87",x"e0",x"c0",x"02"),
  1561 => (x"b7",x"c4",x"49",x"73"),
  1562 => (x"e4",x"c1",x"91",x"29"),
  1563 => (x"4a",x"73",x"81",x"e0"),
  1564 => (x"92",x"c2",x"9a",x"cf"),
  1565 => (x"30",x"72",x"48",x"c1"),
  1566 => (x"ba",x"ff",x"4a",x"70"),
  1567 => (x"98",x"69",x"48",x"72"),
  1568 => (x"87",x"db",x"79",x"70"),
  1569 => (x"b7",x"c4",x"49",x"73"),
  1570 => (x"e4",x"c1",x"91",x"29"),
  1571 => (x"4a",x"73",x"81",x"e0"),
  1572 => (x"92",x"c2",x"9a",x"cf"),
  1573 => (x"30",x"72",x"48",x"c3"),
  1574 => (x"69",x"48",x"4a",x"70"),
  1575 => (x"c1",x"79",x"70",x"b0"),
  1576 => (x"c0",x"48",x"c4",x"e3"),
  1577 => (x"c0",x"e3",x"c1",x"78"),
  1578 => (x"c2",x"78",x"c0",x"48"),
  1579 => (x"f8",x"49",x"fb",x"de"),
  1580 => (x"4a",x"70",x"87",x"e5"),
  1581 => (x"03",x"aa",x"b7",x"c0"),
  1582 => (x"c0",x"87",x"f3",x"fd"),
  1583 => (x"87",x"e4",x"fc",x"48"),
  1584 => (x"00",x"00",x"00",x"00"),
  1585 => (x"00",x"00",x"00",x"00"),
  1586 => (x"49",x"4a",x"71",x"1e"),
  1587 => (x"26",x"87",x"cc",x"fd"),
  1588 => (x"4a",x"c0",x"1e",x"4f"),
  1589 => (x"91",x"c4",x"49",x"72"),
  1590 => (x"81",x"e0",x"e4",x"c1"),
  1591 => (x"82",x"c1",x"79",x"c0"),
  1592 => (x"04",x"aa",x"b7",x"d0"),
  1593 => (x"4f",x"26",x"87",x"ee"),
  1594 => (x"5c",x"5b",x"5e",x"0e"),
  1595 => (x"4d",x"71",x"0e",x"5d"),
  1596 => (x"75",x"87",x"d4",x"f7"),
  1597 => (x"2a",x"b7",x"c4",x"4a"),
  1598 => (x"e0",x"e4",x"c1",x"92"),
  1599 => (x"cf",x"4c",x"75",x"82"),
  1600 => (x"6a",x"94",x"c2",x"9c"),
  1601 => (x"2b",x"74",x"4b",x"49"),
  1602 => (x"48",x"c2",x"9b",x"c3"),
  1603 => (x"4c",x"70",x"30",x"74"),
  1604 => (x"48",x"74",x"bc",x"ff"),
  1605 => (x"7a",x"70",x"98",x"71"),
  1606 => (x"73",x"87",x"e4",x"f6"),
  1607 => (x"87",x"c0",x"fb",x"48"),
  1608 => (x"00",x"00",x"00",x"00"),
  1609 => (x"00",x"00",x"00",x"00"),
  1610 => (x"00",x"00",x"00",x"00"),
  1611 => (x"00",x"00",x"00",x"00"),
  1612 => (x"00",x"00",x"00",x"00"),
  1613 => (x"00",x"00",x"00",x"00"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"00",x"00",x"00",x"00"),
  1616 => (x"00",x"00",x"00",x"00"),
  1617 => (x"00",x"00",x"00",x"00"),
  1618 => (x"00",x"00",x"00",x"00"),
  1619 => (x"00",x"00",x"00",x"00"),
  1620 => (x"00",x"00",x"00",x"00"),
  1621 => (x"00",x"00",x"00",x"00"),
  1622 => (x"00",x"00",x"00",x"00"),
  1623 => (x"00",x"00",x"00",x"00"),
  1624 => (x"25",x"26",x"1e",x"16"),
  1625 => (x"3e",x"3d",x"36",x"2e"),
  1626 => (x"48",x"d0",x"ff",x"1e"),
  1627 => (x"71",x"78",x"e1",x"c8"),
  1628 => (x"08",x"d4",x"ff",x"48"),
  1629 => (x"48",x"66",x"c4",x"78"),
  1630 => (x"78",x"08",x"d4",x"ff"),
  1631 => (x"71",x"1e",x"4f",x"26"),
  1632 => (x"49",x"66",x"c4",x"4a"),
  1633 => (x"ff",x"49",x"72",x"1e"),
  1634 => (x"d0",x"ff",x"87",x"de"),
  1635 => (x"78",x"e0",x"c0",x"48"),
  1636 => (x"1e",x"4f",x"26",x"26"),
  1637 => (x"b7",x"c2",x"4a",x"71"),
  1638 => (x"87",x"c3",x"03",x"aa"),
  1639 => (x"ce",x"87",x"c2",x"82"),
  1640 => (x"1e",x"66",x"c4",x"82"),
  1641 => (x"d5",x"ff",x"49",x"72"),
  1642 => (x"4f",x"26",x"26",x"87"),
  1643 => (x"4a",x"d4",x"ff",x"1e"),
  1644 => (x"ff",x"7a",x"ff",x"c3"),
  1645 => (x"e1",x"c8",x"48",x"d0"),
  1646 => (x"c2",x"7a",x"de",x"78"),
  1647 => (x"7a",x"bf",x"c5",x"df"),
  1648 => (x"28",x"c8",x"48",x"49"),
  1649 => (x"48",x"71",x"7a",x"70"),
  1650 => (x"7a",x"70",x"28",x"d0"),
  1651 => (x"28",x"d8",x"48",x"71"),
  1652 => (x"d0",x"ff",x"7a",x"70"),
  1653 => (x"78",x"e0",x"c0",x"48"),
  1654 => (x"5e",x"0e",x"4f",x"26"),
  1655 => (x"0e",x"5d",x"5c",x"5b"),
  1656 => (x"df",x"c2",x"4c",x"71"),
  1657 => (x"4b",x"4d",x"bf",x"c5"),
  1658 => (x"66",x"d0",x"2b",x"74"),
  1659 => (x"d4",x"83",x"c1",x"9b"),
  1660 => (x"c2",x"04",x"ab",x"66"),
  1661 => (x"74",x"4b",x"c0",x"87"),
  1662 => (x"49",x"66",x"d0",x"4a"),
  1663 => (x"b9",x"ff",x"31",x"72"),
  1664 => (x"48",x"73",x"99",x"75"),
  1665 => (x"4a",x"70",x"30",x"72"),
  1666 => (x"c2",x"b0",x"71",x"48"),
  1667 => (x"fe",x"58",x"c9",x"df"),
  1668 => (x"4d",x"26",x"87",x"da"),
  1669 => (x"4b",x"26",x"4c",x"26"),
  1670 => (x"ff",x"1e",x"4f",x"26"),
  1671 => (x"c9",x"c8",x"48",x"d0"),
  1672 => (x"ff",x"48",x"71",x"78"),
  1673 => (x"26",x"78",x"08",x"d4"),
  1674 => (x"4a",x"71",x"1e",x"4f"),
  1675 => (x"ff",x"87",x"eb",x"49"),
  1676 => (x"78",x"c8",x"48",x"d0"),
  1677 => (x"73",x"1e",x"4f",x"26"),
  1678 => (x"c2",x"4b",x"71",x"1e"),
  1679 => (x"02",x"bf",x"d5",x"df"),
  1680 => (x"eb",x"c2",x"87",x"c3"),
  1681 => (x"48",x"d0",x"ff",x"87"),
  1682 => (x"73",x"78",x"c9",x"c8"),
  1683 => (x"b1",x"e0",x"c0",x"49"),
  1684 => (x"71",x"48",x"d4",x"ff"),
  1685 => (x"c9",x"df",x"c2",x"78"),
  1686 => (x"c8",x"78",x"c0",x"48"),
  1687 => (x"87",x"c5",x"02",x"66"),
  1688 => (x"c2",x"49",x"ff",x"c3"),
  1689 => (x"c2",x"49",x"c0",x"87"),
  1690 => (x"cc",x"59",x"d1",x"df"),
  1691 => (x"87",x"c6",x"02",x"66"),
  1692 => (x"4a",x"d5",x"d5",x"c5"),
  1693 => (x"ff",x"cf",x"87",x"c4"),
  1694 => (x"df",x"c2",x"4a",x"ff"),
  1695 => (x"df",x"c2",x"5a",x"d5"),
  1696 => (x"78",x"c1",x"48",x"d5"),
  1697 => (x"4d",x"26",x"87",x"c4"),
  1698 => (x"4b",x"26",x"4c",x"26"),
  1699 => (x"5e",x"0e",x"4f",x"26"),
  1700 => (x"0e",x"5d",x"5c",x"5b"),
  1701 => (x"df",x"c2",x"4a",x"71"),
  1702 => (x"72",x"4c",x"bf",x"d1"),
  1703 => (x"87",x"cb",x"02",x"9a"),
  1704 => (x"c1",x"91",x"c8",x"49"),
  1705 => (x"71",x"4b",x"ec",x"e8"),
  1706 => (x"c1",x"87",x"c4",x"83"),
  1707 => (x"c0",x"4b",x"ec",x"ec"),
  1708 => (x"74",x"49",x"13",x"4d"),
  1709 => (x"cd",x"df",x"c2",x"99"),
  1710 => (x"d4",x"ff",x"b9",x"bf"),
  1711 => (x"c1",x"78",x"71",x"48"),
  1712 => (x"c8",x"85",x"2c",x"b7"),
  1713 => (x"e8",x"04",x"ad",x"b7"),
  1714 => (x"c9",x"df",x"c2",x"87"),
  1715 => (x"80",x"c8",x"48",x"bf"),
  1716 => (x"58",x"cd",x"df",x"c2"),
  1717 => (x"1e",x"87",x"ef",x"fe"),
  1718 => (x"4b",x"71",x"1e",x"73"),
  1719 => (x"02",x"9a",x"4a",x"13"),
  1720 => (x"49",x"72",x"87",x"cb"),
  1721 => (x"13",x"87",x"e7",x"fe"),
  1722 => (x"f5",x"05",x"9a",x"4a"),
  1723 => (x"87",x"da",x"fe",x"87"),
  1724 => (x"c9",x"df",x"c2",x"1e"),
  1725 => (x"df",x"c2",x"49",x"bf"),
  1726 => (x"a1",x"c1",x"48",x"c9"),
  1727 => (x"b7",x"c0",x"c4",x"78"),
  1728 => (x"87",x"db",x"03",x"a9"),
  1729 => (x"c2",x"48",x"d4",x"ff"),
  1730 => (x"78",x"bf",x"cd",x"df"),
  1731 => (x"bf",x"c9",x"df",x"c2"),
  1732 => (x"c9",x"df",x"c2",x"49"),
  1733 => (x"78",x"a1",x"c1",x"48"),
  1734 => (x"a9",x"b7",x"c0",x"c4"),
  1735 => (x"ff",x"87",x"e5",x"04"),
  1736 => (x"78",x"c8",x"48",x"d0"),
  1737 => (x"48",x"d5",x"df",x"c2"),
  1738 => (x"4f",x"26",x"78",x"c0"),
  1739 => (x"00",x"00",x"00",x"00"),
  1740 => (x"00",x"00",x"00",x"00"),
  1741 => (x"5f",x"00",x"00",x"00"),
  1742 => (x"00",x"00",x"00",x"5f"),
  1743 => (x"00",x"03",x"03",x"00"),
  1744 => (x"00",x"00",x"03",x"03"),
  1745 => (x"14",x"7f",x"7f",x"14"),
  1746 => (x"00",x"14",x"7f",x"7f"),
  1747 => (x"6b",x"2e",x"24",x"00"),
  1748 => (x"00",x"12",x"3a",x"6b"),
  1749 => (x"18",x"36",x"6a",x"4c"),
  1750 => (x"00",x"32",x"56",x"6c"),
  1751 => (x"59",x"4f",x"7e",x"30"),
  1752 => (x"40",x"68",x"3a",x"77"),
  1753 => (x"07",x"04",x"00",x"00"),
  1754 => (x"00",x"00",x"00",x"03"),
  1755 => (x"3e",x"1c",x"00",x"00"),
  1756 => (x"00",x"00",x"41",x"63"),
  1757 => (x"63",x"41",x"00",x"00"),
  1758 => (x"00",x"00",x"1c",x"3e"),
  1759 => (x"1c",x"3e",x"2a",x"08"),
  1760 => (x"08",x"2a",x"3e",x"1c"),
  1761 => (x"3e",x"08",x"08",x"00"),
  1762 => (x"00",x"08",x"08",x"3e"),
  1763 => (x"e0",x"80",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"60"),
  1765 => (x"08",x"08",x"08",x"00"),
  1766 => (x"00",x"08",x"08",x"08"),
  1767 => (x"60",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"60"),
  1769 => (x"18",x"30",x"60",x"40"),
  1770 => (x"01",x"03",x"06",x"0c"),
  1771 => (x"59",x"7f",x"3e",x"00"),
  1772 => (x"00",x"3e",x"7f",x"4d"),
  1773 => (x"7f",x"06",x"04",x"00"),
  1774 => (x"00",x"00",x"00",x"7f"),
  1775 => (x"71",x"63",x"42",x"00"),
  1776 => (x"00",x"46",x"4f",x"59"),
  1777 => (x"49",x"63",x"22",x"00"),
  1778 => (x"00",x"36",x"7f",x"49"),
  1779 => (x"13",x"16",x"1c",x"18"),
  1780 => (x"00",x"10",x"7f",x"7f"),
  1781 => (x"45",x"67",x"27",x"00"),
  1782 => (x"00",x"39",x"7d",x"45"),
  1783 => (x"4b",x"7e",x"3c",x"00"),
  1784 => (x"00",x"30",x"79",x"49"),
  1785 => (x"71",x"01",x"01",x"00"),
  1786 => (x"00",x"07",x"0f",x"79"),
  1787 => (x"49",x"7f",x"36",x"00"),
  1788 => (x"00",x"36",x"7f",x"49"),
  1789 => (x"49",x"4f",x"06",x"00"),
  1790 => (x"00",x"1e",x"3f",x"69"),
  1791 => (x"66",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"66"),
  1793 => (x"e6",x"80",x"00",x"00"),
  1794 => (x"00",x"00",x"00",x"66"),
  1795 => (x"14",x"08",x"08",x"00"),
  1796 => (x"00",x"22",x"22",x"14"),
  1797 => (x"14",x"14",x"14",x"00"),
  1798 => (x"00",x"14",x"14",x"14"),
  1799 => (x"14",x"22",x"22",x"00"),
  1800 => (x"00",x"08",x"08",x"14"),
  1801 => (x"51",x"03",x"02",x"00"),
  1802 => (x"00",x"06",x"0f",x"59"),
  1803 => (x"5d",x"41",x"7f",x"3e"),
  1804 => (x"00",x"1e",x"1f",x"55"),
  1805 => (x"09",x"7f",x"7e",x"00"),
  1806 => (x"00",x"7e",x"7f",x"09"),
  1807 => (x"49",x"7f",x"7f",x"00"),
  1808 => (x"00",x"36",x"7f",x"49"),
  1809 => (x"63",x"3e",x"1c",x"00"),
  1810 => (x"00",x"41",x"41",x"41"),
  1811 => (x"41",x"7f",x"7f",x"00"),
  1812 => (x"00",x"1c",x"3e",x"63"),
  1813 => (x"49",x"7f",x"7f",x"00"),
  1814 => (x"00",x"41",x"41",x"49"),
  1815 => (x"09",x"7f",x"7f",x"00"),
  1816 => (x"00",x"01",x"01",x"09"),
  1817 => (x"41",x"7f",x"3e",x"00"),
  1818 => (x"00",x"7a",x"7b",x"49"),
  1819 => (x"08",x"7f",x"7f",x"00"),
  1820 => (x"00",x"7f",x"7f",x"08"),
  1821 => (x"7f",x"41",x"00",x"00"),
  1822 => (x"00",x"00",x"41",x"7f"),
  1823 => (x"40",x"60",x"20",x"00"),
  1824 => (x"00",x"3f",x"7f",x"40"),
  1825 => (x"1c",x"08",x"7f",x"7f"),
  1826 => (x"00",x"41",x"63",x"36"),
  1827 => (x"40",x"7f",x"7f",x"00"),
  1828 => (x"00",x"40",x"40",x"40"),
  1829 => (x"0c",x"06",x"7f",x"7f"),
  1830 => (x"00",x"7f",x"7f",x"06"),
  1831 => (x"0c",x"06",x"7f",x"7f"),
  1832 => (x"00",x"7f",x"7f",x"18"),
  1833 => (x"41",x"7f",x"3e",x"00"),
  1834 => (x"00",x"3e",x"7f",x"41"),
  1835 => (x"09",x"7f",x"7f",x"00"),
  1836 => (x"00",x"06",x"0f",x"09"),
  1837 => (x"61",x"41",x"7f",x"3e"),
  1838 => (x"00",x"40",x"7e",x"7f"),
  1839 => (x"09",x"7f",x"7f",x"00"),
  1840 => (x"00",x"66",x"7f",x"19"),
  1841 => (x"4d",x"6f",x"26",x"00"),
  1842 => (x"00",x"32",x"7b",x"59"),
  1843 => (x"7f",x"01",x"01",x"00"),
  1844 => (x"00",x"01",x"01",x"7f"),
  1845 => (x"40",x"7f",x"3f",x"00"),
  1846 => (x"00",x"3f",x"7f",x"40"),
  1847 => (x"70",x"3f",x"0f",x"00"),
  1848 => (x"00",x"0f",x"3f",x"70"),
  1849 => (x"18",x"30",x"7f",x"7f"),
  1850 => (x"00",x"7f",x"7f",x"30"),
  1851 => (x"1c",x"36",x"63",x"41"),
  1852 => (x"41",x"63",x"36",x"1c"),
  1853 => (x"7c",x"06",x"03",x"01"),
  1854 => (x"01",x"03",x"06",x"7c"),
  1855 => (x"4d",x"59",x"71",x"61"),
  1856 => (x"00",x"41",x"43",x"47"),
  1857 => (x"7f",x"7f",x"00",x"00"),
  1858 => (x"00",x"00",x"41",x"41"),
  1859 => (x"0c",x"06",x"03",x"01"),
  1860 => (x"40",x"60",x"30",x"18"),
  1861 => (x"41",x"41",x"00",x"00"),
  1862 => (x"00",x"00",x"7f",x"7f"),
  1863 => (x"03",x"06",x"0c",x"08"),
  1864 => (x"00",x"08",x"0c",x"06"),
  1865 => (x"80",x"80",x"80",x"80"),
  1866 => (x"00",x"80",x"80",x"80"),
  1867 => (x"03",x"00",x"00",x"00"),
  1868 => (x"00",x"00",x"04",x"07"),
  1869 => (x"54",x"74",x"20",x"00"),
  1870 => (x"00",x"78",x"7c",x"54"),
  1871 => (x"44",x"7f",x"7f",x"00"),
  1872 => (x"00",x"38",x"7c",x"44"),
  1873 => (x"44",x"7c",x"38",x"00"),
  1874 => (x"00",x"00",x"44",x"44"),
  1875 => (x"44",x"7c",x"38",x"00"),
  1876 => (x"00",x"7f",x"7f",x"44"),
  1877 => (x"54",x"7c",x"38",x"00"),
  1878 => (x"00",x"18",x"5c",x"54"),
  1879 => (x"7f",x"7e",x"04",x"00"),
  1880 => (x"00",x"00",x"05",x"05"),
  1881 => (x"a4",x"bc",x"18",x"00"),
  1882 => (x"00",x"7c",x"fc",x"a4"),
  1883 => (x"04",x"7f",x"7f",x"00"),
  1884 => (x"00",x"78",x"7c",x"04"),
  1885 => (x"3d",x"00",x"00",x"00"),
  1886 => (x"00",x"00",x"40",x"7d"),
  1887 => (x"80",x"80",x"80",x"00"),
  1888 => (x"00",x"00",x"7d",x"fd"),
  1889 => (x"10",x"7f",x"7f",x"00"),
  1890 => (x"00",x"44",x"6c",x"38"),
  1891 => (x"3f",x"00",x"00",x"00"),
  1892 => (x"00",x"00",x"40",x"7f"),
  1893 => (x"18",x"0c",x"7c",x"7c"),
  1894 => (x"00",x"78",x"7c",x"0c"),
  1895 => (x"04",x"7c",x"7c",x"00"),
  1896 => (x"00",x"78",x"7c",x"04"),
  1897 => (x"44",x"7c",x"38",x"00"),
  1898 => (x"00",x"38",x"7c",x"44"),
  1899 => (x"24",x"fc",x"fc",x"00"),
  1900 => (x"00",x"18",x"3c",x"24"),
  1901 => (x"24",x"3c",x"18",x"00"),
  1902 => (x"00",x"fc",x"fc",x"24"),
  1903 => (x"04",x"7c",x"7c",x"00"),
  1904 => (x"00",x"08",x"0c",x"04"),
  1905 => (x"54",x"5c",x"48",x"00"),
  1906 => (x"00",x"20",x"74",x"54"),
  1907 => (x"7f",x"3f",x"04",x"00"),
  1908 => (x"00",x"00",x"44",x"44"),
  1909 => (x"40",x"7c",x"3c",x"00"),
  1910 => (x"00",x"7c",x"7c",x"40"),
  1911 => (x"60",x"3c",x"1c",x"00"),
  1912 => (x"00",x"1c",x"3c",x"60"),
  1913 => (x"30",x"60",x"7c",x"3c"),
  1914 => (x"00",x"3c",x"7c",x"60"),
  1915 => (x"10",x"38",x"6c",x"44"),
  1916 => (x"00",x"44",x"6c",x"38"),
  1917 => (x"e0",x"bc",x"1c",x"00"),
  1918 => (x"00",x"1c",x"3c",x"60"),
  1919 => (x"74",x"64",x"44",x"00"),
  1920 => (x"00",x"44",x"4c",x"5c"),
  1921 => (x"3e",x"08",x"08",x"00"),
  1922 => (x"00",x"41",x"41",x"77"),
  1923 => (x"7f",x"00",x"00",x"00"),
  1924 => (x"00",x"00",x"00",x"7f"),
  1925 => (x"77",x"41",x"41",x"00"),
  1926 => (x"00",x"08",x"08",x"3e"),
  1927 => (x"03",x"01",x"01",x"02"),
  1928 => (x"00",x"01",x"02",x"02"),
  1929 => (x"7f",x"7f",x"7f",x"7f"),
  1930 => (x"00",x"7f",x"7f",x"7f"),
  1931 => (x"1c",x"1c",x"08",x"08"),
  1932 => (x"7f",x"7f",x"3e",x"3e"),
  1933 => (x"3e",x"3e",x"7f",x"7f"),
  1934 => (x"08",x"08",x"1c",x"1c"),
  1935 => (x"7c",x"18",x"10",x"00"),
  1936 => (x"00",x"10",x"18",x"7c"),
  1937 => (x"7c",x"30",x"10",x"00"),
  1938 => (x"00",x"10",x"30",x"7c"),
  1939 => (x"60",x"60",x"30",x"10"),
  1940 => (x"00",x"06",x"1e",x"78"),
  1941 => (x"18",x"3c",x"66",x"42"),
  1942 => (x"00",x"42",x"66",x"3c"),
  1943 => (x"c2",x"6a",x"38",x"78"),
  1944 => (x"00",x"38",x"6c",x"c6"),
  1945 => (x"60",x"00",x"00",x"60"),
  1946 => (x"00",x"60",x"00",x"00"),
  1947 => (x"5c",x"5b",x"5e",x"0e"),
  1948 => (x"71",x"1e",x"0e",x"5d"),
  1949 => (x"e6",x"df",x"c2",x"4c"),
  1950 => (x"4b",x"c0",x"4d",x"bf"),
  1951 => (x"ab",x"74",x"1e",x"c0"),
  1952 => (x"c4",x"87",x"c7",x"02"),
  1953 => (x"78",x"c0",x"48",x"a6"),
  1954 => (x"a6",x"c4",x"87",x"c5"),
  1955 => (x"c4",x"78",x"c1",x"48"),
  1956 => (x"49",x"73",x"1e",x"66"),
  1957 => (x"c8",x"87",x"df",x"ee"),
  1958 => (x"49",x"e0",x"c0",x"86"),
  1959 => (x"c4",x"87",x"ef",x"ef"),
  1960 => (x"49",x"6a",x"4a",x"a5"),
  1961 => (x"f1",x"87",x"f0",x"f0"),
  1962 => (x"85",x"cb",x"87",x"c6"),
  1963 => (x"b7",x"c8",x"83",x"c1"),
  1964 => (x"c7",x"ff",x"04",x"ab"),
  1965 => (x"4d",x"26",x"26",x"87"),
  1966 => (x"4b",x"26",x"4c",x"26"),
  1967 => (x"71",x"1e",x"4f",x"26"),
  1968 => (x"ea",x"df",x"c2",x"4a"),
  1969 => (x"ea",x"df",x"c2",x"5a"),
  1970 => (x"49",x"78",x"c7",x"48"),
  1971 => (x"26",x"87",x"dd",x"fe"),
  1972 => (x"1e",x"73",x"1e",x"4f"),
  1973 => (x"b7",x"c0",x"4a",x"71"),
  1974 => (x"87",x"d3",x"03",x"aa"),
  1975 => (x"bf",x"e1",x"c8",x"c2"),
  1976 => (x"c1",x"87",x"c4",x"05"),
  1977 => (x"c0",x"87",x"c2",x"4b"),
  1978 => (x"e5",x"c8",x"c2",x"4b"),
  1979 => (x"c2",x"87",x"c4",x"5b"),
  1980 => (x"c2",x"5a",x"e5",x"c8"),
  1981 => (x"4a",x"bf",x"e1",x"c8"),
  1982 => (x"c0",x"c1",x"9a",x"c1"),
  1983 => (x"e8",x"ec",x"49",x"a2"),
  1984 => (x"c2",x"48",x"fc",x"87"),
  1985 => (x"78",x"bf",x"e1",x"c8"),
  1986 => (x"1e",x"87",x"ef",x"fe"),
  1987 => (x"66",x"c4",x"4a",x"71"),
  1988 => (x"e9",x"49",x"72",x"1e"),
  1989 => (x"26",x"26",x"87",x"fd"),
  1990 => (x"c8",x"c2",x"1e",x"4f"),
  1991 => (x"e6",x"49",x"bf",x"e1"),
  1992 => (x"df",x"c2",x"87",x"e6"),
  1993 => (x"bf",x"e8",x"48",x"de"),
  1994 => (x"da",x"df",x"c2",x"78"),
  1995 => (x"78",x"bf",x"ec",x"48"),
  1996 => (x"bf",x"de",x"df",x"c2"),
  1997 => (x"ff",x"c3",x"49",x"4a"),
  1998 => (x"2a",x"b7",x"c8",x"99"),
  1999 => (x"b0",x"71",x"48",x"72"),
  2000 => (x"58",x"e6",x"df",x"c2"),
  2001 => (x"5e",x"0e",x"4f",x"26"),
  2002 => (x"0e",x"5d",x"5c",x"5b"),
  2003 => (x"c8",x"ff",x"4b",x"71"),
  2004 => (x"d9",x"df",x"c2",x"87"),
  2005 => (x"73",x"50",x"c0",x"48"),
  2006 => (x"87",x"cc",x"e6",x"49"),
  2007 => (x"c2",x"4c",x"49",x"70"),
  2008 => (x"49",x"ee",x"cb",x"9c"),
  2009 => (x"70",x"87",x"c2",x"cb"),
  2010 => (x"df",x"c2",x"4d",x"49"),
  2011 => (x"05",x"bf",x"97",x"d9"),
  2012 => (x"d0",x"87",x"e2",x"c1"),
  2013 => (x"df",x"c2",x"49",x"66"),
  2014 => (x"05",x"99",x"bf",x"e2"),
  2015 => (x"66",x"d4",x"87",x"d6"),
  2016 => (x"da",x"df",x"c2",x"49"),
  2017 => (x"cb",x"05",x"99",x"bf"),
  2018 => (x"e5",x"49",x"73",x"87"),
  2019 => (x"98",x"70",x"87",x"da"),
  2020 => (x"87",x"c1",x"c1",x"02"),
  2021 => (x"c0",x"fe",x"4c",x"c1"),
  2022 => (x"ca",x"49",x"75",x"87"),
  2023 => (x"98",x"70",x"87",x"d7"),
  2024 => (x"c2",x"87",x"c6",x"02"),
  2025 => (x"c1",x"48",x"d9",x"df"),
  2026 => (x"d9",x"df",x"c2",x"50"),
  2027 => (x"c0",x"05",x"bf",x"97"),
  2028 => (x"df",x"c2",x"87",x"e3"),
  2029 => (x"d0",x"49",x"bf",x"e2"),
  2030 => (x"ff",x"05",x"99",x"66"),
  2031 => (x"df",x"c2",x"87",x"d6"),
  2032 => (x"d4",x"49",x"bf",x"da"),
  2033 => (x"ff",x"05",x"99",x"66"),
  2034 => (x"49",x"73",x"87",x"ca"),
  2035 => (x"70",x"87",x"d9",x"e4"),
  2036 => (x"ff",x"fe",x"05",x"98"),
  2037 => (x"fb",x"48",x"74",x"87"),
  2038 => (x"5e",x"0e",x"87",x"dc"),
  2039 => (x"0e",x"5d",x"5c",x"5b"),
  2040 => (x"4d",x"c0",x"86",x"f4"),
  2041 => (x"7e",x"bf",x"ec",x"4c"),
  2042 => (x"c2",x"48",x"a6",x"c4"),
  2043 => (x"78",x"bf",x"e6",x"df"),
  2044 => (x"1e",x"c0",x"1e",x"c1"),
  2045 => (x"cd",x"fd",x"49",x"c7"),
  2046 => (x"70",x"86",x"c8",x"87"),
  2047 => (x"87",x"cd",x"02",x"98"),
  2048 => (x"cc",x"fb",x"49",x"ff"),
  2049 => (x"49",x"da",x"c1",x"87"),
  2050 => (x"c1",x"87",x"dd",x"e3"),
  2051 => (x"d9",x"df",x"c2",x"4d"),
  2052 => (x"c3",x"02",x"bf",x"97"),
  2053 => (x"87",x"f3",x"cc",x"87"),
  2054 => (x"bf",x"de",x"df",x"c2"),
  2055 => (x"e1",x"c8",x"c2",x"4b"),
  2056 => (x"e9",x"c0",x"05",x"bf"),
  2057 => (x"49",x"fd",x"c3",x"87"),
  2058 => (x"c3",x"87",x"fd",x"e2"),
  2059 => (x"f7",x"e2",x"49",x"fa"),
  2060 => (x"c3",x"49",x"73",x"87"),
  2061 => (x"1e",x"71",x"99",x"ff"),
  2062 => (x"ce",x"fb",x"49",x"c0"),
  2063 => (x"c8",x"49",x"73",x"87"),
  2064 => (x"1e",x"71",x"29",x"b7"),
  2065 => (x"c2",x"fb",x"49",x"c1"),
  2066 => (x"c5",x"86",x"c8",x"87"),
  2067 => (x"df",x"c2",x"87",x"f9"),
  2068 => (x"9b",x"4b",x"bf",x"e2"),
  2069 => (x"c2",x"87",x"dd",x"02"),
  2070 => (x"49",x"bf",x"dd",x"c8"),
  2071 => (x"70",x"87",x"d6",x"c7"),
  2072 => (x"87",x"c4",x"05",x"98"),
  2073 => (x"87",x"d2",x"4b",x"c0"),
  2074 => (x"c6",x"49",x"e0",x"c2"),
  2075 => (x"c8",x"c2",x"87",x"fb"),
  2076 => (x"87",x"c6",x"58",x"e1"),
  2077 => (x"48",x"dd",x"c8",x"c2"),
  2078 => (x"49",x"73",x"78",x"c0"),
  2079 => (x"cd",x"05",x"99",x"c2"),
  2080 => (x"49",x"eb",x"c3",x"87"),
  2081 => (x"70",x"87",x"e1",x"e1"),
  2082 => (x"02",x"99",x"c2",x"49"),
  2083 => (x"4c",x"fb",x"87",x"c2"),
  2084 => (x"99",x"c1",x"49",x"73"),
  2085 => (x"c3",x"87",x"cd",x"05"),
  2086 => (x"cb",x"e1",x"49",x"f4"),
  2087 => (x"c2",x"49",x"70",x"87"),
  2088 => (x"87",x"c2",x"02",x"99"),
  2089 => (x"49",x"73",x"4c",x"fa"),
  2090 => (x"cd",x"05",x"99",x"c8"),
  2091 => (x"49",x"f5",x"c3",x"87"),
  2092 => (x"70",x"87",x"f5",x"e0"),
  2093 => (x"02",x"99",x"c2",x"49"),
  2094 => (x"df",x"c2",x"87",x"d4"),
  2095 => (x"c9",x"02",x"bf",x"ea"),
  2096 => (x"88",x"c1",x"48",x"87"),
  2097 => (x"58",x"ee",x"df",x"c2"),
  2098 => (x"4c",x"ff",x"87",x"c2"),
  2099 => (x"49",x"73",x"4d",x"c1"),
  2100 => (x"cd",x"05",x"99",x"c4"),
  2101 => (x"49",x"f2",x"c3",x"87"),
  2102 => (x"70",x"87",x"cd",x"e0"),
  2103 => (x"02",x"99",x"c2",x"49"),
  2104 => (x"df",x"c2",x"87",x"db"),
  2105 => (x"48",x"7e",x"bf",x"ea"),
  2106 => (x"03",x"a8",x"b7",x"c7"),
  2107 => (x"48",x"6e",x"87",x"cb"),
  2108 => (x"df",x"c2",x"80",x"c1"),
  2109 => (x"c2",x"c0",x"58",x"ee"),
  2110 => (x"c1",x"4c",x"fe",x"87"),
  2111 => (x"49",x"fd",x"c3",x"4d"),
  2112 => (x"87",x"e4",x"df",x"ff"),
  2113 => (x"99",x"c2",x"49",x"70"),
  2114 => (x"c2",x"87",x"d5",x"02"),
  2115 => (x"02",x"bf",x"ea",x"df"),
  2116 => (x"c2",x"87",x"c9",x"c0"),
  2117 => (x"c0",x"48",x"ea",x"df"),
  2118 => (x"87",x"c2",x"c0",x"78"),
  2119 => (x"4d",x"c1",x"4c",x"fd"),
  2120 => (x"ff",x"49",x"fa",x"c3"),
  2121 => (x"70",x"87",x"c1",x"df"),
  2122 => (x"02",x"99",x"c2",x"49"),
  2123 => (x"df",x"c2",x"87",x"d9"),
  2124 => (x"c7",x"48",x"bf",x"ea"),
  2125 => (x"c0",x"03",x"a8",x"b7"),
  2126 => (x"df",x"c2",x"87",x"c9"),
  2127 => (x"78",x"c7",x"48",x"ea"),
  2128 => (x"fc",x"87",x"c2",x"c0"),
  2129 => (x"c0",x"4d",x"c1",x"4c"),
  2130 => (x"c0",x"03",x"ac",x"b7"),
  2131 => (x"66",x"c4",x"87",x"d1"),
  2132 => (x"82",x"d8",x"c1",x"4a"),
  2133 => (x"c6",x"c0",x"02",x"6a"),
  2134 => (x"74",x"4b",x"6a",x"87"),
  2135 => (x"c0",x"0f",x"73",x"49"),
  2136 => (x"1e",x"f0",x"c3",x"1e"),
  2137 => (x"f7",x"49",x"da",x"c1"),
  2138 => (x"86",x"c8",x"87",x"dc"),
  2139 => (x"c0",x"02",x"98",x"70"),
  2140 => (x"a6",x"c8",x"87",x"e2"),
  2141 => (x"ea",x"df",x"c2",x"48"),
  2142 => (x"66",x"c8",x"78",x"bf"),
  2143 => (x"c4",x"91",x"cb",x"49"),
  2144 => (x"80",x"71",x"48",x"66"),
  2145 => (x"bf",x"6e",x"7e",x"70"),
  2146 => (x"87",x"c8",x"c0",x"02"),
  2147 => (x"c8",x"4b",x"bf",x"6e"),
  2148 => (x"0f",x"73",x"49",x"66"),
  2149 => (x"c0",x"02",x"9d",x"75"),
  2150 => (x"df",x"c2",x"87",x"c8"),
  2151 => (x"f3",x"49",x"bf",x"ea"),
  2152 => (x"c8",x"c2",x"87",x"ca"),
  2153 => (x"c0",x"02",x"bf",x"e5"),
  2154 => (x"c2",x"49",x"87",x"dd"),
  2155 => (x"98",x"70",x"87",x"c7"),
  2156 => (x"87",x"d3",x"c0",x"02"),
  2157 => (x"bf",x"ea",x"df",x"c2"),
  2158 => (x"87",x"f0",x"f2",x"49"),
  2159 => (x"d0",x"f4",x"49",x"c0"),
  2160 => (x"e5",x"c8",x"c2",x"87"),
  2161 => (x"f4",x"78",x"c0",x"48"),
  2162 => (x"87",x"ea",x"f3",x"8e"),
  2163 => (x"5c",x"5b",x"5e",x"0e"),
  2164 => (x"71",x"1e",x"0e",x"5d"),
  2165 => (x"e6",x"df",x"c2",x"4c"),
  2166 => (x"cd",x"c1",x"49",x"bf"),
  2167 => (x"d1",x"c1",x"4d",x"a1"),
  2168 => (x"74",x"7e",x"69",x"81"),
  2169 => (x"87",x"cf",x"02",x"9c"),
  2170 => (x"74",x"4b",x"a5",x"c4"),
  2171 => (x"e6",x"df",x"c2",x"7b"),
  2172 => (x"c9",x"f3",x"49",x"bf"),
  2173 => (x"74",x"7b",x"6e",x"87"),
  2174 => (x"87",x"c4",x"05",x"9c"),
  2175 => (x"87",x"c2",x"4b",x"c0"),
  2176 => (x"49",x"73",x"4b",x"c1"),
  2177 => (x"d4",x"87",x"ca",x"f3"),
  2178 => (x"87",x"c7",x"02",x"66"),
  2179 => (x"70",x"87",x"da",x"49"),
  2180 => (x"c0",x"87",x"c2",x"4a"),
  2181 => (x"e9",x"c8",x"c2",x"4a"),
  2182 => (x"d9",x"f2",x"26",x"5a"),
  2183 => (x"00",x"00",x"00",x"87"),
  2184 => (x"00",x"00",x"00",x"00"),
  2185 => (x"00",x"00",x"00",x"00"),
  2186 => (x"4a",x"71",x"1e",x"00"),
  2187 => (x"49",x"bf",x"c8",x"ff"),
  2188 => (x"26",x"48",x"a1",x"72"),
  2189 => (x"c8",x"ff",x"1e",x"4f"),
  2190 => (x"c0",x"fe",x"89",x"bf"),
  2191 => (x"c0",x"c0",x"c0",x"c0"),
  2192 => (x"87",x"c4",x"01",x"a9"),
  2193 => (x"87",x"c2",x"4a",x"c0"),
  2194 => (x"48",x"72",x"4a",x"c1"),
  2195 => (x"5e",x"0e",x"4f",x"26"),
  2196 => (x"0e",x"5d",x"5c",x"5b"),
  2197 => (x"ff",x"7e",x"71",x"1e"),
  2198 => (x"1e",x"6e",x"4b",x"d4"),
  2199 => (x"49",x"ee",x"df",x"c2"),
  2200 => (x"87",x"f1",x"d5",x"fe"),
  2201 => (x"4d",x"70",x"86",x"c4"),
  2202 => (x"c3",x"c3",x"02",x"9d"),
  2203 => (x"f6",x"df",x"c2",x"87"),
  2204 => (x"49",x"6e",x"4c",x"bf"),
  2205 => (x"87",x"e6",x"e7",x"fe"),
  2206 => (x"c8",x"48",x"d0",x"ff"),
  2207 => (x"d6",x"c1",x"78",x"c5"),
  2208 => (x"15",x"4a",x"c0",x"7b"),
  2209 => (x"c0",x"82",x"c1",x"7b"),
  2210 => (x"04",x"aa",x"b7",x"e0"),
  2211 => (x"d0",x"ff",x"87",x"f5"),
  2212 => (x"c8",x"78",x"c4",x"48"),
  2213 => (x"d3",x"c1",x"78",x"c5"),
  2214 => (x"c4",x"7b",x"c1",x"7b"),
  2215 => (x"02",x"9c",x"74",x"78"),
  2216 => (x"c2",x"87",x"fc",x"c1"),
  2217 => (x"c8",x"7e",x"de",x"ce"),
  2218 => (x"c0",x"8c",x"4d",x"c0"),
  2219 => (x"c6",x"03",x"ac",x"b7"),
  2220 => (x"a4",x"c0",x"c8",x"87"),
  2221 => (x"c2",x"4c",x"c0",x"4d"),
  2222 => (x"bf",x"97",x"cf",x"db"),
  2223 => (x"02",x"99",x"d0",x"49"),
  2224 => (x"1e",x"c0",x"87",x"d2"),
  2225 => (x"49",x"ee",x"df",x"c2"),
  2226 => (x"87",x"e5",x"d7",x"fe"),
  2227 => (x"49",x"70",x"86",x"c4"),
  2228 => (x"87",x"ef",x"c0",x"4a"),
  2229 => (x"1e",x"de",x"ce",x"c2"),
  2230 => (x"49",x"ee",x"df",x"c2"),
  2231 => (x"87",x"d1",x"d7",x"fe"),
  2232 => (x"49",x"70",x"86",x"c4"),
  2233 => (x"48",x"d0",x"ff",x"4a"),
  2234 => (x"c1",x"78",x"c5",x"c8"),
  2235 => (x"97",x"6e",x"7b",x"d4"),
  2236 => (x"48",x"6e",x"7b",x"bf"),
  2237 => (x"7e",x"70",x"80",x"c1"),
  2238 => (x"ff",x"05",x"8d",x"c1"),
  2239 => (x"d0",x"ff",x"87",x"f0"),
  2240 => (x"72",x"78",x"c4",x"48"),
  2241 => (x"87",x"c5",x"05",x"9a"),
  2242 => (x"e5",x"c0",x"48",x"c0"),
  2243 => (x"c2",x"1e",x"c1",x"87"),
  2244 => (x"fe",x"49",x"ee",x"df"),
  2245 => (x"c4",x"87",x"f9",x"d4"),
  2246 => (x"05",x"9c",x"74",x"86"),
  2247 => (x"ff",x"87",x"c4",x"fe"),
  2248 => (x"c5",x"c8",x"48",x"d0"),
  2249 => (x"7b",x"d3",x"c1",x"78"),
  2250 => (x"78",x"c4",x"7b",x"c0"),
  2251 => (x"87",x"c2",x"48",x"c1"),
  2252 => (x"26",x"26",x"48",x"c0"),
  2253 => (x"26",x"4c",x"26",x"4d"),
  2254 => (x"1e",x"4f",x"26",x"4b"),
  2255 => (x"66",x"c4",x"4a",x"71"),
  2256 => (x"72",x"87",x"c5",x"05"),
  2257 => (x"87",x"c6",x"fc",x"49"),
  2258 => (x"1e",x"00",x"4f",x"26"),
  2259 => (x"bf",x"f4",x"cd",x"c2"),
  2260 => (x"c2",x"b9",x"c1",x"49"),
  2261 => (x"ff",x"59",x"f8",x"cd"),
  2262 => (x"ff",x"c3",x"48",x"d4"),
  2263 => (x"48",x"d0",x"ff",x"78"),
  2264 => (x"ff",x"78",x"e1",x"c8"),
  2265 => (x"78",x"c1",x"48",x"d4"),
  2266 => (x"78",x"71",x"31",x"c4"),
  2267 => (x"c0",x"48",x"d0",x"ff"),
  2268 => (x"4f",x"26",x"78",x"e0"),
  2269 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

